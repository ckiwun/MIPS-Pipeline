
module DataMemory_test_1 ( clk, rst, stall, EX_WB, EX_MEM, EX_ALUresult, 
        EX_RegisterRd, MEMWriteData, WB, MemoryData, ALUresult, RegisterRd, 
        read_MemoryData, test_si, test_so, test_se );
  input [1:0] EX_WB;
  input [2:0] EX_MEM;
  input [31:0] EX_ALUresult;
  input [4:0] EX_RegisterRd;
  input [31:0] MEMWriteData;
  output [1:0] WB;
  output [31:0] MemoryData;
  output [31:0] ALUresult;
  output [4:0] RegisterRd;
  input [31:0] read_MemoryData;
  input clk, rst, stall, test_si, test_se;
  output test_so;
  wire   n169, n170, n171, n172, n173, n174, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n1, n34,
         n35, n36, n37, n38, n39, n40, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n156, n157, n158, n159, n160, n161;

  CLKBUFX2 U2 ( .A(stall), .Y(n40) );
  MX2XL U3 ( .A(EX_RegisterRd[0]), .B(RegisterRd[0]), .S0(n145), .Y(n107) );
  MX2XL U4 ( .A(EX_RegisterRd[1]), .B(RegisterRd[1]), .S0(n145), .Y(n108) );
  MX2XL U5 ( .A(EX_RegisterRd[3]), .B(RegisterRd[3]), .S0(n145), .Y(n110) );
  MX2XL U6 ( .A(EX_RegisterRd[2]), .B(RegisterRd[2]), .S0(n145), .Y(n109) );
  MX2XL U7 ( .A(EX_RegisterRd[4]), .B(RegisterRd[4]), .S0(n145), .Y(n111) );
  MX2XL U8 ( .A(EX_WB[1]), .B(WB[1]), .S0(n144), .Y(n106) );
  INVX3 U9 ( .A(n40), .Y(n36) );
  INVX3 U10 ( .A(n40), .Y(n37) );
  INVX3 U11 ( .A(n40), .Y(n38) );
  INVX3 U12 ( .A(n144), .Y(n35) );
  INVX3 U13 ( .A(n144), .Y(n34) );
  INVX3 U14 ( .A(n40), .Y(n39) );
  CLKBUFX3 U15 ( .A(n1), .Y(n145) );
  CLKBUFX3 U16 ( .A(n1), .Y(n144) );
  CLKBUFX3 U17 ( .A(n153), .Y(n147) );
  CLKBUFX3 U18 ( .A(n153), .Y(n148) );
  CLKBUFX3 U19 ( .A(n146), .Y(n149) );
  CLKBUFX3 U20 ( .A(n153), .Y(n150) );
  CLKBUFX3 U21 ( .A(n146), .Y(n151) );
  CLKBUFX3 U22 ( .A(n146), .Y(n152) );
  CLKBUFX3 U23 ( .A(stall), .Y(n1) );
  CLKBUFX3 U24 ( .A(n146), .Y(n153) );
  CLKBUFX3 U25 ( .A(rst), .Y(n146) );
  OAI2BB2XL U26 ( .B0(n41), .B1(n34), .A0N(EX_ALUresult[0]), .A1N(n37), .Y(
        n112) );
  OAI2BB2XL U27 ( .B0(n42), .B1(n35), .A0N(EX_ALUresult[1]), .A1N(n36), .Y(
        n113) );
  OAI2BB2XL U28 ( .B0(n43), .B1(n35), .A0N(EX_ALUresult[2]), .A1N(n36), .Y(
        n114) );
  OAI2BB2XL U29 ( .B0(n44), .B1(n34), .A0N(EX_ALUresult[3]), .A1N(n37), .Y(
        n115) );
  OAI2BB2XL U30 ( .B0(n45), .B1(n35), .A0N(EX_ALUresult[4]), .A1N(n37), .Y(
        n116) );
  OAI2BB2XL U31 ( .B0(n46), .B1(n34), .A0N(EX_ALUresult[5]), .A1N(n37), .Y(
        n117) );
  OAI2BB2XL U32 ( .B0(n47), .B1(n36), .A0N(EX_ALUresult[6]), .A1N(n38), .Y(
        n118) );
  OAI2BB2XL U33 ( .B0(n48), .B1(n34), .A0N(EX_ALUresult[7]), .A1N(n38), .Y(
        n119) );
  OAI2BB2XL U34 ( .B0(n49), .B1(n34), .A0N(EX_ALUresult[8]), .A1N(n37), .Y(
        n120) );
  OAI2BB2XL U35 ( .B0(n50), .B1(n34), .A0N(EX_ALUresult[9]), .A1N(n37), .Y(
        n121) );
  OAI2BB2XL U36 ( .B0(n51), .B1(n34), .A0N(EX_ALUresult[10]), .A1N(n37), .Y(
        n122) );
  OAI2BB2XL U37 ( .B0(n52), .B1(n34), .A0N(EX_ALUresult[11]), .A1N(n37), .Y(
        n123) );
  OAI2BB2XL U38 ( .B0(n53), .B1(n34), .A0N(EX_ALUresult[12]), .A1N(n38), .Y(
        n124) );
  OAI2BB2XL U39 ( .B0(n54), .B1(n34), .A0N(EX_ALUresult[13]), .A1N(n37), .Y(
        n125) );
  OAI2BB2XL U40 ( .B0(n55), .B1(n34), .A0N(EX_ALUresult[14]), .A1N(n38), .Y(
        n126) );
  OAI2BB2XL U41 ( .B0(n56), .B1(n34), .A0N(EX_ALUresult[15]), .A1N(n38), .Y(
        n127) );
  OAI2BB2XL U42 ( .B0(n57), .B1(n34), .A0N(EX_ALUresult[16]), .A1N(n38), .Y(
        n128) );
  OAI2BB2XL U43 ( .B0(n58), .B1(n34), .A0N(EX_ALUresult[17]), .A1N(n38), .Y(
        n129) );
  OAI2BB2XL U44 ( .B0(n59), .B1(n34), .A0N(EX_ALUresult[18]), .A1N(n38), .Y(
        n130) );
  OAI2BB2XL U45 ( .B0(n60), .B1(n39), .A0N(EX_ALUresult[19]), .A1N(n38), .Y(
        n131) );
  OAI2BB2XL U46 ( .B0(n61), .B1(n39), .A0N(EX_ALUresult[20]), .A1N(n38), .Y(
        n132) );
  OAI2BB2XL U47 ( .B0(n62), .B1(n39), .A0N(EX_ALUresult[21]), .A1N(n39), .Y(
        n133) );
  OAI2BB2XL U48 ( .B0(n63), .B1(n39), .A0N(EX_ALUresult[22]), .A1N(n38), .Y(
        n134) );
  OAI2BB2XL U49 ( .B0(n64), .B1(n35), .A0N(EX_ALUresult[23]), .A1N(n38), .Y(
        n135) );
  OAI2BB2XL U50 ( .B0(n65), .B1(n34), .A0N(EX_ALUresult[24]), .A1N(n39), .Y(
        n136) );
  OAI2BB2XL U51 ( .B0(n66), .B1(n34), .A0N(EX_ALUresult[25]), .A1N(n39), .Y(
        n137) );
  OAI2BB2XL U52 ( .B0(n67), .B1(n34), .A0N(EX_ALUresult[26]), .A1N(n39), .Y(
        n138) );
  OAI2BB2XL U53 ( .B0(n68), .B1(n39), .A0N(EX_ALUresult[27]), .A1N(n39), .Y(
        n139) );
  OAI2BB2XL U54 ( .B0(n69), .B1(n36), .A0N(EX_ALUresult[28]), .A1N(n39), .Y(
        n140) );
  OAI2BB2XL U55 ( .B0(n70), .B1(n35), .A0N(EX_ALUresult[29]), .A1N(n39), .Y(
        n141) );
  OAI2BB2XL U56 ( .B0(n71), .B1(n38), .A0N(EX_ALUresult[30]), .A1N(n39), .Y(
        n142) );
  OAI2BB2XL U57 ( .B0(n72), .B1(n39), .A0N(EX_ALUresult[31]), .A1N(n39), .Y(
        n143) );
  OAI2BB2XL U58 ( .B0(n2), .B1(n36), .A0N(read_MemoryData[0]), .A1N(n39), .Y(
        n73) );
  OAI2BB2XL U59 ( .B0(n3), .B1(n35), .A0N(read_MemoryData[1]), .A1N(n39), .Y(
        n74) );
  OAI2BB2XL U60 ( .B0(n4), .B1(n36), .A0N(read_MemoryData[2]), .A1N(n39), .Y(
        n75) );
  OAI2BB2XL U61 ( .B0(n5), .B1(n35), .A0N(read_MemoryData[3]), .A1N(n39), .Y(
        n76) );
  OAI2BB2XL U62 ( .B0(n6), .B1(n35), .A0N(read_MemoryData[4]), .A1N(n38), .Y(
        n77) );
  OAI2BB2XL U63 ( .B0(n7), .B1(n36), .A0N(read_MemoryData[5]), .A1N(n38), .Y(
        n78) );
  OAI2BB2XL U64 ( .B0(n8), .B1(n36), .A0N(read_MemoryData[6]), .A1N(n38), .Y(
        n79) );
  OAI2BB2XL U65 ( .B0(n9), .B1(n35), .A0N(read_MemoryData[7]), .A1N(n38), .Y(
        n80) );
  OAI2BB2XL U66 ( .B0(n10), .B1(n35), .A0N(read_MemoryData[8]), .A1N(n38), .Y(
        n81) );
  OAI2BB2XL U67 ( .B0(n11), .B1(n35), .A0N(read_MemoryData[9]), .A1N(n38), .Y(
        n82) );
  OAI2BB2XL U68 ( .B0(n12), .B1(n36), .A0N(read_MemoryData[10]), .A1N(n37), 
        .Y(n83) );
  OAI2BB2XL U69 ( .B0(n13), .B1(n35), .A0N(read_MemoryData[11]), .A1N(n37), 
        .Y(n84) );
  OAI2BB2XL U70 ( .B0(n14), .B1(n35), .A0N(read_MemoryData[12]), .A1N(n37), 
        .Y(n85) );
  OAI2BB2XL U71 ( .B0(n15), .B1(n35), .A0N(read_MemoryData[13]), .A1N(n37), 
        .Y(n86) );
  OAI2BB2XL U72 ( .B0(n16), .B1(n35), .A0N(read_MemoryData[14]), .A1N(n38), 
        .Y(n87) );
  OAI2BB2XL U73 ( .B0(n17), .B1(n35), .A0N(read_MemoryData[15]), .A1N(n37), 
        .Y(n88) );
  OAI2BB2XL U74 ( .B0(n18), .B1(n39), .A0N(read_MemoryData[16]), .A1N(n36), 
        .Y(n89) );
  OAI2BB2XL U75 ( .B0(n19), .B1(n37), .A0N(read_MemoryData[17]), .A1N(n37), 
        .Y(n90) );
  OAI2BB2XL U76 ( .B0(n20), .B1(n35), .A0N(read_MemoryData[18]), .A1N(n36), 
        .Y(n91) );
  OAI2BB2XL U77 ( .B0(n21), .B1(n35), .A0N(read_MemoryData[19]), .A1N(n37), 
        .Y(n92) );
  OAI2BB2XL U78 ( .B0(n22), .B1(n34), .A0N(read_MemoryData[20]), .A1N(n36), 
        .Y(n93) );
  OAI2BB2XL U79 ( .B0(n23), .B1(n38), .A0N(read_MemoryData[21]), .A1N(n37), 
        .Y(n94) );
  OAI2BB2XL U80 ( .B0(n24), .B1(n36), .A0N(read_MemoryData[22]), .A1N(n36), 
        .Y(n95) );
  OAI2BB2XL U81 ( .B0(n25), .B1(n39), .A0N(read_MemoryData[23]), .A1N(n36), 
        .Y(n96) );
  OAI2BB2XL U82 ( .B0(n26), .B1(n37), .A0N(read_MemoryData[24]), .A1N(n36), 
        .Y(n97) );
  OAI2BB2XL U83 ( .B0(n27), .B1(n35), .A0N(read_MemoryData[25]), .A1N(n37), 
        .Y(n98) );
  OAI2BB2XL U84 ( .B0(n28), .B1(n34), .A0N(read_MemoryData[26]), .A1N(n36), 
        .Y(n99) );
  OAI2BB2XL U85 ( .B0(n29), .B1(n34), .A0N(read_MemoryData[27]), .A1N(n36), 
        .Y(n100) );
  OAI2BB2XL U86 ( .B0(n30), .B1(n35), .A0N(read_MemoryData[28]), .A1N(n36), 
        .Y(n101) );
  OAI2BB2XL U87 ( .B0(n31), .B1(n35), .A0N(read_MemoryData[29]), .A1N(n37), 
        .Y(n102) );
  OAI2BB2XL U88 ( .B0(n32), .B1(n37), .A0N(read_MemoryData[30]), .A1N(n36), 
        .Y(n103) );
  OAI2BB2XL U89 ( .B0(n33), .B1(n38), .A0N(read_MemoryData[31]), .A1N(n36), 
        .Y(n104) );
  CLKMX2X2 U90 ( .A(EX_WB[0]), .B(WB[0]), .S0(n144), .Y(n105) );
  SDFFRXL \MemoryData_reg[31]  ( .D(n104), .SI(n32), .SE(test_se), .CK(clk), 
        .RN(n149), .Q(MemoryData[31]), .QN(n33) );
  SDFFRXL \MemoryData_reg[30]  ( .D(n103), .SI(n31), .SE(test_se), .CK(clk), 
        .RN(n149), .Q(MemoryData[30]), .QN(n32) );
  SDFFRXL \MemoryData_reg[29]  ( .D(n102), .SI(n30), .SE(test_se), .CK(clk), 
        .RN(n149), .Q(MemoryData[29]), .QN(n31) );
  SDFFRXL \MemoryData_reg[28]  ( .D(n101), .SI(n29), .SE(test_se), .CK(clk), 
        .RN(n149), .Q(MemoryData[28]), .QN(n30) );
  SDFFRXL \MemoryData_reg[27]  ( .D(n100), .SI(n28), .SE(test_se), .CK(clk), 
        .RN(n149), .Q(MemoryData[27]), .QN(n29) );
  SDFFRXL \MemoryData_reg[26]  ( .D(n99), .SI(n27), .SE(test_se), .CK(clk), 
        .RN(n149), .Q(MemoryData[26]), .QN(n28) );
  SDFFRXL \MemoryData_reg[25]  ( .D(n98), .SI(n26), .SE(test_se), .CK(clk), 
        .RN(n149), .Q(MemoryData[25]), .QN(n27) );
  SDFFRXL \MemoryData_reg[24]  ( .D(n97), .SI(n25), .SE(test_se), .CK(clk), 
        .RN(n149), .Q(MemoryData[24]), .QN(n26) );
  SDFFRXL \MemoryData_reg[23]  ( .D(n96), .SI(n24), .SE(test_se), .CK(clk), 
        .RN(n148), .Q(MemoryData[23]), .QN(n25) );
  SDFFRXL \MemoryData_reg[22]  ( .D(n95), .SI(n23), .SE(test_se), .CK(clk), 
        .RN(n148), .Q(MemoryData[22]), .QN(n24) );
  SDFFRXL \MemoryData_reg[21]  ( .D(n94), .SI(n22), .SE(test_se), .CK(clk), 
        .RN(n148), .Q(MemoryData[21]), .QN(n23) );
  SDFFRXL \MemoryData_reg[20]  ( .D(n93), .SI(n21), .SE(test_se), .CK(clk), 
        .RN(n148), .Q(MemoryData[20]), .QN(n22) );
  SDFFRXL \MemoryData_reg[19]  ( .D(n92), .SI(n20), .SE(test_se), .CK(clk), 
        .RN(n148), .Q(MemoryData[19]), .QN(n21) );
  SDFFRXL \MemoryData_reg[18]  ( .D(n91), .SI(n19), .SE(test_se), .CK(clk), 
        .RN(n148), .Q(MemoryData[18]), .QN(n20) );
  SDFFRXL \MemoryData_reg[17]  ( .D(n90), .SI(n18), .SE(test_se), .CK(clk), 
        .RN(n148), .Q(MemoryData[17]), .QN(n19) );
  SDFFRXL \MemoryData_reg[16]  ( .D(n89), .SI(n17), .SE(test_se), .CK(clk), 
        .RN(n148), .Q(MemoryData[16]), .QN(n18) );
  SDFFRXL \MemoryData_reg[15]  ( .D(n88), .SI(n16), .SE(test_se), .CK(clk), 
        .RN(n148), .Q(MemoryData[15]), .QN(n17) );
  SDFFRXL \MemoryData_reg[14]  ( .D(n87), .SI(n15), .SE(test_se), .CK(clk), 
        .RN(n148), .Q(MemoryData[14]), .QN(n16) );
  SDFFRXL \MemoryData_reg[13]  ( .D(n86), .SI(n14), .SE(test_se), .CK(clk), 
        .RN(n148), .Q(MemoryData[13]), .QN(n15) );
  SDFFRXL \MemoryData_reg[12]  ( .D(n85), .SI(n13), .SE(test_se), .CK(clk), 
        .RN(n148), .Q(MemoryData[12]), .QN(n14) );
  SDFFRXL \MemoryData_reg[11]  ( .D(n84), .SI(n12), .SE(test_se), .CK(clk), 
        .RN(n147), .Q(MemoryData[11]), .QN(n13) );
  SDFFRXL \MemoryData_reg[10]  ( .D(n83), .SI(n11), .SE(test_se), .CK(clk), 
        .RN(n147), .Q(MemoryData[10]), .QN(n12) );
  SDFFRXL \MemoryData_reg[9]  ( .D(n82), .SI(n10), .SE(test_se), .CK(clk), 
        .RN(n147), .Q(MemoryData[9]), .QN(n11) );
  SDFFRXL \MemoryData_reg[8]  ( .D(n81), .SI(n9), .SE(test_se), .CK(clk), .RN(
        n147), .Q(MemoryData[8]), .QN(n10) );
  SDFFRXL \MemoryData_reg[7]  ( .D(n80), .SI(n8), .SE(test_se), .CK(clk), .RN(
        n147), .Q(MemoryData[7]), .QN(n9) );
  SDFFRXL \MemoryData_reg[6]  ( .D(n79), .SI(n7), .SE(test_se), .CK(clk), .RN(
        n147), .Q(MemoryData[6]), .QN(n8) );
  SDFFRXL \MemoryData_reg[5]  ( .D(n78), .SI(n6), .SE(test_se), .CK(clk), .RN(
        n147), .Q(MemoryData[5]), .QN(n7) );
  SDFFRXL \MemoryData_reg[4]  ( .D(n77), .SI(n5), .SE(test_se), .CK(clk), .RN(
        n147), .Q(MemoryData[4]), .QN(n6) );
  SDFFRXL \MemoryData_reg[3]  ( .D(n76), .SI(n4), .SE(test_se), .CK(clk), .RN(
        n147), .Q(MemoryData[3]), .QN(n5) );
  SDFFRXL \MemoryData_reg[2]  ( .D(n75), .SI(n3), .SE(test_se), .CK(clk), .RN(
        n147), .Q(MemoryData[2]), .QN(n4) );
  SDFFRXL \MemoryData_reg[1]  ( .D(n74), .SI(n2), .SE(test_se), .CK(clk), .RN(
        n147), .Q(MemoryData[1]), .QN(n3) );
  SDFFRXL \MemoryData_reg[0]  ( .D(n73), .SI(n72), .SE(test_se), .CK(clk), 
        .RN(n147), .Q(MemoryData[0]), .QN(n2) );
  SDFFRXL \ALUresult_reg[31]  ( .D(n143), .SI(n71), .SE(test_se), .CK(clk), 
        .RN(n152), .Q(ALUresult[31]), .QN(n72) );
  SDFFRXL \ALUresult_reg[30]  ( .D(n142), .SI(n70), .SE(test_se), .CK(clk), 
        .RN(n152), .Q(ALUresult[30]), .QN(n71) );
  SDFFRXL \ALUresult_reg[29]  ( .D(n141), .SI(n69), .SE(test_se), .CK(clk), 
        .RN(n152), .Q(ALUresult[29]), .QN(n70) );
  SDFFRXL \ALUresult_reg[28]  ( .D(n140), .SI(n68), .SE(test_se), .CK(clk), 
        .RN(n152), .Q(ALUresult[28]), .QN(n69) );
  SDFFRXL \ALUresult_reg[27]  ( .D(n139), .SI(n67), .SE(test_se), .CK(clk), 
        .RN(n152), .Q(ALUresult[27]), .QN(n68) );
  SDFFRXL \ALUresult_reg[26]  ( .D(n138), .SI(n66), .SE(test_se), .CK(clk), 
        .RN(n152), .Q(ALUresult[26]), .QN(n67) );
  SDFFRXL \ALUresult_reg[25]  ( .D(n137), .SI(n65), .SE(test_se), .CK(clk), 
        .RN(n152), .Q(ALUresult[25]), .QN(n66) );
  SDFFRXL \ALUresult_reg[24]  ( .D(n136), .SI(n64), .SE(test_se), .CK(clk), 
        .RN(n152), .Q(ALUresult[24]), .QN(n65) );
  SDFFRXL \ALUresult_reg[23]  ( .D(n135), .SI(n63), .SE(test_se), .CK(clk), 
        .RN(n152), .Q(ALUresult[23]), .QN(n64) );
  SDFFRXL \ALUresult_reg[22]  ( .D(n134), .SI(n62), .SE(test_se), .CK(clk), 
        .RN(n152), .Q(ALUresult[22]), .QN(n63) );
  SDFFRXL \ALUresult_reg[21]  ( .D(n133), .SI(n61), .SE(test_se), .CK(clk), 
        .RN(n152), .Q(ALUresult[21]), .QN(n62) );
  SDFFRXL \ALUresult_reg[20]  ( .D(n132), .SI(n60), .SE(test_se), .CK(clk), 
        .RN(n151), .Q(ALUresult[20]), .QN(n61) );
  SDFFRXL \ALUresult_reg[19]  ( .D(n131), .SI(n59), .SE(test_se), .CK(clk), 
        .RN(n151), .Q(ALUresult[19]), .QN(n60) );
  SDFFRXL \ALUresult_reg[18]  ( .D(n130), .SI(n58), .SE(test_se), .CK(clk), 
        .RN(n151), .Q(ALUresult[18]), .QN(n59) );
  SDFFRXL \ALUresult_reg[17]  ( .D(n129), .SI(n57), .SE(test_se), .CK(clk), 
        .RN(n151), .Q(ALUresult[17]), .QN(n58) );
  SDFFRXL \ALUresult_reg[16]  ( .D(n128), .SI(n56), .SE(test_se), .CK(clk), 
        .RN(n151), .Q(ALUresult[16]), .QN(n57) );
  SDFFRXL \ALUresult_reg[15]  ( .D(n127), .SI(n55), .SE(test_se), .CK(clk), 
        .RN(n151), .Q(ALUresult[15]), .QN(n56) );
  SDFFRXL \ALUresult_reg[14]  ( .D(n126), .SI(n54), .SE(test_se), .CK(clk), 
        .RN(n151), .Q(ALUresult[14]), .QN(n55) );
  SDFFRXL \ALUresult_reg[13]  ( .D(n125), .SI(n53), .SE(test_se), .CK(clk), 
        .RN(n151), .Q(ALUresult[13]), .QN(n54) );
  SDFFRXL \ALUresult_reg[12]  ( .D(n124), .SI(n52), .SE(test_se), .CK(clk), 
        .RN(n151), .Q(ALUresult[12]), .QN(n53) );
  SDFFRXL \ALUresult_reg[11]  ( .D(n123), .SI(n51), .SE(test_se), .CK(clk), 
        .RN(n151), .Q(ALUresult[11]), .QN(n52) );
  SDFFRXL \ALUresult_reg[10]  ( .D(n122), .SI(n50), .SE(test_se), .CK(clk), 
        .RN(n151), .Q(ALUresult[10]), .QN(n51) );
  SDFFRXL \ALUresult_reg[9]  ( .D(n121), .SI(n49), .SE(test_se), .CK(clk), 
        .RN(n151), .Q(ALUresult[9]), .QN(n50) );
  SDFFRXL \ALUresult_reg[8]  ( .D(n120), .SI(n48), .SE(test_se), .CK(clk), 
        .RN(n150), .Q(ALUresult[8]), .QN(n49) );
  SDFFRXL \ALUresult_reg[7]  ( .D(n119), .SI(n47), .SE(test_se), .CK(clk), 
        .RN(n150), .Q(ALUresult[7]), .QN(n48) );
  SDFFRXL \ALUresult_reg[6]  ( .D(n118), .SI(n46), .SE(test_se), .CK(clk), 
        .RN(n150), .Q(ALUresult[6]), .QN(n47) );
  SDFFRXL \ALUresult_reg[5]  ( .D(n117), .SI(n45), .SE(test_se), .CK(clk), 
        .RN(n150), .Q(ALUresult[5]), .QN(n46) );
  SDFFRXL \ALUresult_reg[4]  ( .D(n116), .SI(n44), .SE(test_se), .CK(clk), 
        .RN(n150), .Q(ALUresult[4]), .QN(n45) );
  SDFFRXL \ALUresult_reg[3]  ( .D(n115), .SI(n43), .SE(test_se), .CK(clk), 
        .RN(n150), .Q(ALUresult[3]), .QN(n44) );
  SDFFRXL \ALUresult_reg[2]  ( .D(n114), .SI(n42), .SE(test_se), .CK(clk), 
        .RN(n150), .Q(ALUresult[2]), .QN(n43) );
  SDFFRXL \ALUresult_reg[1]  ( .D(n113), .SI(n41), .SE(test_se), .CK(clk), 
        .RN(n150), .Q(ALUresult[1]), .QN(n42) );
  SDFFRXL \ALUresult_reg[0]  ( .D(n112), .SI(test_si), .SE(test_se), .CK(clk), 
        .RN(n150), .Q(ALUresult[0]), .QN(n41) );
  SDFFRXL \WB_reg[1]  ( .D(n106), .SI(n158), .SE(test_se), .CK(clk), .RN(n149), 
        .Q(n169), .QN(test_so) );
  SDFFRXL \RegisterRd_reg[1]  ( .D(n108), .SI(n156), .SE(test_se), .CK(clk), 
        .RN(n149), .Q(n173), .QN(n161) );
  SDFFRXL \RegisterRd_reg[2]  ( .D(n109), .SI(n161), .SE(test_se), .CK(clk), 
        .RN(n150), .Q(n172), .QN(n160) );
  SDFFRXL \RegisterRd_reg[3]  ( .D(n110), .SI(n160), .SE(test_se), .CK(clk), 
        .RN(n150), .Q(n171), .QN(n159) );
  SDFFRXL \WB_reg[0]  ( .D(n105), .SI(n157), .SE(test_se), .CK(clk), .RN(rst), 
        .Q(WB[0]), .QN(n158) );
  SDFFRXL \RegisterRd_reg[4]  ( .D(n111), .SI(n159), .SE(test_se), .CK(clk), 
        .RN(n150), .Q(n170), .QN(n157) );
  SDFFRXL \RegisterRd_reg[0]  ( .D(n107), .SI(n33), .SE(test_se), .CK(clk), 
        .RN(n149), .Q(n174), .QN(n156) );
  CLKBUFX2 U1 ( .A(n170), .Y(RegisterRd[4]) );
  CLKBUFX2 U91 ( .A(n169), .Y(WB[1]) );
  CLKBUFX2 U92 ( .A(n172), .Y(RegisterRd[2]) );
  CLKBUFX2 U93 ( .A(n171), .Y(RegisterRd[3]) );
  CLKBUFX2 U94 ( .A(n174), .Y(RegisterRd[0]) );
  CLKBUFX2 U95 ( .A(n173), .Y(RegisterRd[1]) );
endmodule


module Execution_DW_cmp_0 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375;

  CLKINVX1 U654 ( .A(B[27]), .Y(n1283) );
  CLKINVX1 U655 ( .A(B[31]), .Y(n1278) );
  CLKINVX1 U656 ( .A(B[30]), .Y(n1279) );
  OAI21XL U657 ( .A0(n1332), .A1(n1333), .B0(n1334), .Y(n1317) );
  AOI32XL U658 ( .A0(B[2]), .A1(n1311), .A2(n1374), .B0(n1310), .B1(B[3]), .Y(
        n1372) );
  OAI211X1 U659 ( .A0(B[12]), .A1(n1301), .B0(n1360), .C0(n1358), .Y(n1353) );
  INVXL U660 ( .A(A[13]), .Y(n1300) );
  NAND2BXL U661 ( .AN(B[13]), .B(A[13]), .Y(n1360) );
  AOI32XL U662 ( .A0(B[12]), .A1(n1301), .A2(n1360), .B0(n1300), .B1(B[13]), 
        .Y(n1359) );
  CLKINVX1 U663 ( .A(B[1]), .Y(n1312) );
  AOI21XL U664 ( .A0(n1284), .A1(A[26]), .B0(n1344), .Y(n1342) );
  OAI211X1 U665 ( .A0(B[8]), .A1(n1305), .B0(n1351), .C0(n1352), .Y(n1350) );
  AOI32XL U666 ( .A0(B[8]), .A1(n1305), .A2(n1351), .B0(n1304), .B1(B[9]), .Y(
        n1363) );
  AND2XL U667 ( .A(A[15]), .B(n1297), .Y(n1361) );
  OAI22XL U668 ( .A0(n1340), .A1(n1341), .B0(n1342), .B1(n1340), .Y(n1333) );
  OAI22XL U669 ( .A0(n1335), .A1(n1280), .B0(n1336), .B1(n1335), .Y(n1334) );
  OAI32XL U670 ( .A0(n1289), .A1(A[22]), .A2(n1325), .B0(A[23]), .B1(n1288), 
        .Y(n1321) );
  OAI32XL U671 ( .A0(n1307), .A1(A[6]), .A2(n1369), .B0(A[7]), .B1(n1306), .Y(
        n1365) );
  OAI32XL U672 ( .A0(n1293), .A1(A[18]), .A2(n1330), .B0(A[19]), .B1(n1292), 
        .Y(n1326) );
  AOI211XL U673 ( .A0(n1291), .A1(A[20]), .B0(n1324), .C0(n1323), .Y(n1331) );
  INVXL U674 ( .A(A[11]), .Y(n1302) );
  AOI21XL U675 ( .A0(n1307), .A1(A[6]), .B0(n1369), .Y(n1367) );
  AOI21XL U676 ( .A0(n1293), .A1(A[18]), .B0(n1330), .Y(n1327) );
  OAI32XL U677 ( .A0(n1291), .A1(A[20]), .A2(n1324), .B0(A[21]), .B1(n1290), 
        .Y(n1322) );
  OAI32XL U678 ( .A0(n1286), .A1(A[24]), .A2(n1343), .B0(A[25]), .B1(n1285), 
        .Y(n1341) );
  OAI211XL U679 ( .A0(B[16]), .A1(n1296), .B0(n1329), .C0(n1346), .Y(n1314) );
  NAND3XL U680 ( .A(n1367), .B(n1370), .C(n1371), .Y(n1347) );
  NAND2BXL U681 ( .AN(B[11]), .B(A[11]), .Y(n1364) );
  INVXL U682 ( .A(A[29]), .Y(n1281) );
  AND2XL U683 ( .A(A[25]), .B(n1285), .Y(n1343) );
  AND2XL U684 ( .A(A[21]), .B(n1290), .Y(n1324) );
  AND2XL U685 ( .A(A[27]), .B(n1283), .Y(n1344) );
  AND2XL U686 ( .A(A[19]), .B(n1292), .Y(n1330) );
  AND2X2 U687 ( .A(A[31]), .B(n1278), .Y(n1339) );
  AND2XL U688 ( .A(A[7]), .B(n1306), .Y(n1369) );
  AO21XL U689 ( .A0(n1289), .A1(A[22]), .B0(n1325), .Y(n1323) );
  AND2XL U690 ( .A(A[23]), .B(n1288), .Y(n1325) );
  INVXL U691 ( .A(B[26]), .Y(n1284) );
  INVXL U692 ( .A(B[24]), .Y(n1286) );
  INVXL U693 ( .A(B[25]), .Y(n1285) );
  INVXL U694 ( .A(B[23]), .Y(n1288) );
  INVXL U695 ( .A(B[19]), .Y(n1292) );
  INVXL U696 ( .A(B[21]), .Y(n1290) );
  INVXL U697 ( .A(B[0]), .Y(n1313) );
  INVXL U698 ( .A(A[3]), .Y(n1310) );
  NOR2BXL U699 ( .AN(A[5]), .B(B[5]), .Y(n1368) );
  NAND2BXL U700 ( .AN(B[17]), .B(A[17]), .Y(n1329) );
  NAND2BXL U701 ( .AN(B[9]), .B(A[9]), .Y(n1351) );
  NAND2BXL U702 ( .AN(B[3]), .B(A[3]), .Y(n1374) );
  INVXL U703 ( .A(B[20]), .Y(n1291) );
  INVXL U704 ( .A(B[18]), .Y(n1293) );
  INVXL U705 ( .A(B[22]), .Y(n1289) );
  INVXL U706 ( .A(A[16]), .Y(n1296) );
  OAI2BB1X1 U707 ( .A0N(n1331), .A1N(n1277), .B0(n1320), .Y(n1318) );
  OA22X1 U708 ( .A0(n1326), .A1(n1294), .B0(n1327), .B1(n1326), .Y(n1277) );
  CLKINVX1 U709 ( .A(n1323), .Y(n1287) );
  INVXL U710 ( .A(B[14]), .Y(n1298) );
  INVXL U711 ( .A(B[15]), .Y(n1297) );
  CLKINVX1 U712 ( .A(n1359), .Y(n1299) );
  INVXL U713 ( .A(B[5]), .Y(n1308) );
  INVXL U714 ( .A(B[6]), .Y(n1307) );
  INVXL U715 ( .A(B[7]), .Y(n1306) );
  INVXL U716 ( .A(B[4]), .Y(n1309) );
  INVXL U717 ( .A(A[12]), .Y(n1301) );
  INVXL U718 ( .A(A[8]), .Y(n1305) );
  CLKINVX1 U719 ( .A(A[28]), .Y(n1282) );
  INVXL U720 ( .A(A[10]), .Y(n1303) );
  INVXL U721 ( .A(A[2]), .Y(n1311) );
  INVXL U722 ( .A(A[9]), .Y(n1304) );
  CLKINVX1 U723 ( .A(n1328), .Y(n1294) );
  INVXL U724 ( .A(A[17]), .Y(n1295) );
  CLKINVX1 U725 ( .A(n1337), .Y(n1280) );
  OAI21XL U726 ( .A0(n1314), .A1(n1315), .B0(n1316), .Y(GE_LT_GT_LE) );
  OAI22XL U727 ( .A0(n1317), .A1(n1318), .B0(n1319), .B1(n1317), .Y(n1316) );
  OAI22XL U728 ( .A0(n1321), .A1(n1322), .B0(n1287), .B1(n1321), .Y(n1320) );
  AOI32X1 U729 ( .A0(B[16]), .A1(n1296), .A2(n1329), .B0(n1295), .B1(B[17]), 
        .Y(n1328) );
  AOI32X1 U730 ( .A0(B[28]), .A1(n1282), .A2(n1338), .B0(n1281), .B1(B[29]), 
        .Y(n1337) );
  OAI32X1 U731 ( .A0(n1279), .A1(A[30]), .A2(n1339), .B0(A[31]), .B1(n1278), 
        .Y(n1335) );
  OAI32X1 U732 ( .A0(n1284), .A1(A[26]), .A2(n1344), .B0(A[27]), .B1(n1283), 
        .Y(n1340) );
  NAND3X1 U733 ( .A(n1319), .B(n1331), .C(n1327), .Y(n1315) );
  AOI211X1 U734 ( .A0(n1286), .A1(A[24]), .B0(n1343), .C0(n1345), .Y(n1319) );
  NAND2BX1 U735 ( .AN(n1332), .B(n1342), .Y(n1345) );
  OAI211X1 U736 ( .A0(B[28]), .A1(n1282), .B0(n1338), .C0(n1336), .Y(n1332) );
  AOI21X1 U737 ( .A0(n1279), .A1(A[30]), .B0(n1339), .Y(n1336) );
  NAND2BX1 U738 ( .AN(B[29]), .B(A[29]), .Y(n1338) );
  AOI32X1 U739 ( .A0(n1347), .A1(n1348), .A2(n1349), .B0(n1349), .B1(n1350), 
        .Y(n1346) );
  NOR2X1 U740 ( .A(n1353), .B(n1354), .Y(n1352) );
  OA21XL U741 ( .A0(n1353), .A1(n1355), .B0(n1356), .Y(n1349) );
  OAI22XL U742 ( .A0(n1357), .A1(n1299), .B0(n1358), .B1(n1357), .Y(n1356) );
  OAI32X1 U743 ( .A0(n1298), .A1(A[14]), .A2(n1361), .B0(A[15]), .B1(n1297), 
        .Y(n1357) );
  AO22X1 U744 ( .A0(n1362), .A1(n1363), .B0(n1354), .B1(n1362), .Y(n1355) );
  OAI21XL U745 ( .A0(B[10]), .A1(n1303), .B0(n1364), .Y(n1354) );
  AOI32X1 U746 ( .A0(B[10]), .A1(n1303), .A2(n1364), .B0(n1302), .B1(B[11]), 
        .Y(n1362) );
  AOI21X1 U747 ( .A0(n1298), .A1(A[14]), .B0(n1361), .Y(n1358) );
  OAI22XL U748 ( .A0(n1365), .A1(n1366), .B0(n1367), .B1(n1365), .Y(n1348) );
  OAI32X1 U749 ( .A0(n1309), .A1(A[4]), .A2(n1368), .B0(A[5]), .B1(n1308), .Y(
        n1366) );
  AOI221XL U750 ( .A0(n1372), .A1(n1373), .B0(A[4]), .B1(n1309), .C0(n1368), 
        .Y(n1371) );
  OAI21XL U751 ( .A0(B[2]), .A1(n1311), .B0(n1374), .Y(n1373) );
  OAI211X1 U752 ( .A0(A[1]), .A1(n1312), .B0(n1375), .C0(n1372), .Y(n1370) );
  AO22X1 U753 ( .A0(n1313), .A1(A[0]), .B0(n1312), .B1(A[1]), .Y(n1375) );
endmodule


module Execution_DW_rightsh_0 ( A, DATA_TC, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC;
  wire   n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365;

  NOR2BX1 U179 ( .AN(n323), .B(n230), .Y(n310) );
  MXI3X1 U180 ( .A(n284), .B(n248), .C(n285), .S0(n233), .S1(n237), .Y(B[3])
         );
  MXI3X1 U181 ( .A(n273), .B(n309), .C(n292), .S0(n233), .S1(n236), .Y(B[14])
         );
  MXI3X1 U182 ( .A(n283), .B(n313), .C(n301), .S0(n233), .S1(n236), .Y(B[12])
         );
  MXI3X1 U183 ( .A(n258), .B(n259), .C(n260), .S0(n233), .S1(n236), .Y(B[9])
         );
  MXI2XL U184 ( .A(n329), .B(n330), .S0(n231), .Y(n307) );
  MX2XL U185 ( .A(A[13]), .B(A[14]), .S0(n226), .Y(n347) );
  NAND2XL U186 ( .A(n305), .B(n234), .Y(n263) );
  INVXL U187 ( .A(n332), .Y(n249) );
  CLKMX2X2 U188 ( .A(n323), .B(n324), .S0(n231), .Y(n304) );
  NOR2X1 U189 ( .A(n237), .B(n275), .Y(B[21]) );
  MXI3XL U190 ( .A(n268), .B(n307), .C(n291), .S0(n233), .S1(n236), .Y(B[15])
         );
  MXI3XL U191 ( .A(n278), .B(n311), .C(n300), .S0(n233), .S1(n236), .Y(B[13])
         );
  CLKINVX1 U192 ( .A(n271), .Y(n253) );
  NAND2XL U193 ( .A(n320), .B(n234), .Y(n302) );
  NAND2XL U194 ( .A(n322), .B(n234), .Y(n303) );
  NAND2XL U195 ( .A(n306), .B(n234), .Y(n291) );
  NOR2XL U196 ( .A(n237), .B(n270), .Y(B[22]) );
  INVX1 U197 ( .A(n286), .Y(n248) );
  MXI2XL U198 ( .A(A[5]), .B(A[6]), .S0(SH[0]), .Y(n288) );
  MXI2XL U199 ( .A(A[3]), .B(A[4]), .S0(SH[0]), .Y(n287) );
  NOR2BXL U200 ( .AN(A[31]), .B(n226), .Y(n338) );
  MX2XL U201 ( .A(A[0]), .B(A[1]), .S0(n226), .Y(n365) );
  MX2XL U202 ( .A(A[15]), .B(A[16]), .S0(n226), .Y(n346) );
  MX2XL U203 ( .A(A[28]), .B(A[29]), .S0(n226), .Y(n353) );
  MX2XL U204 ( .A(A[26]), .B(A[27]), .S0(n226), .Y(n354) );
  MX2XL U205 ( .A(A[24]), .B(A[25]), .S0(n226), .Y(n358) );
  MX2XL U206 ( .A(A[25]), .B(A[26]), .S0(n226), .Y(n343) );
  MX2XL U207 ( .A(A[22]), .B(A[23]), .S0(n225), .Y(n359) );
  MX2XL U208 ( .A(A[23]), .B(A[24]), .S0(n226), .Y(n340) );
  MX2XL U209 ( .A(A[21]), .B(A[22]), .S0(n226), .Y(n341) );
  MX2XL U210 ( .A(A[18]), .B(A[19]), .S0(n225), .Y(n357) );
  MX2XL U211 ( .A(A[20]), .B(A[21]), .S0(n225), .Y(n356) );
  MX2XL U212 ( .A(A[19]), .B(A[20]), .S0(n226), .Y(n344) );
  MX2XL U213 ( .A(A[7]), .B(A[8]), .S0(n226), .Y(n289) );
  MX2XL U214 ( .A(A[11]), .B(A[12]), .S0(n226), .Y(n318) );
  MX2XL U215 ( .A(A[9]), .B(A[10]), .S0(n225), .Y(n290) );
  MX2XL U216 ( .A(A[8]), .B(A[9]), .S0(n225), .Y(n299) );
  MX2XL U217 ( .A(A[12]), .B(A[13]), .S0(n225), .Y(n361) );
  MX2XL U218 ( .A(A[10]), .B(A[11]), .S0(n225), .Y(n360) );
  MX2XL U219 ( .A(A[16]), .B(A[17]), .S0(n225), .Y(n362) );
  MX2XL U220 ( .A(A[14]), .B(A[15]), .S0(n225), .Y(n363) );
  MX2XL U221 ( .A(A[27]), .B(A[28]), .S0(n226), .Y(n342) );
  MX2XL U222 ( .A(A[6]), .B(A[7]), .S0(n225), .Y(n298) );
  MX2XL U223 ( .A(A[29]), .B(A[30]), .S0(n226), .Y(n339) );
  MX2XL U224 ( .A(A[17]), .B(A[18]), .S0(n226), .Y(n345) );
  MX2XL U225 ( .A(A[4]), .B(A[5]), .S0(n225), .Y(n297) );
  MX2XL U226 ( .A(A[30]), .B(A[31]), .S0(n225), .Y(n355) );
  MX2XL U227 ( .A(A[2]), .B(A[3]), .S0(n225), .Y(n296) );
  CLKINVX1 U228 ( .A(n327), .Y(n239) );
  CLKINVX1 U229 ( .A(n307), .Y(n243) );
  CLKINVX1 U230 ( .A(n309), .Y(n244) );
  CLKINVX1 U231 ( .A(n311), .Y(n245) );
  CLKINVX1 U232 ( .A(n259), .Y(n247) );
  CLKINVX1 U233 ( .A(n313), .Y(n246) );
  CLKINVX1 U234 ( .A(n302), .Y(n238) );
  CLKINVX1 U235 ( .A(n303), .Y(n241) );
  CLKINVX1 U236 ( .A(n263), .Y(n240) );
  INVX3 U237 ( .A(n227), .Y(n228) );
  CLKINVX1 U238 ( .A(n227), .Y(n229) );
  INVX3 U239 ( .A(n230), .Y(n231) );
  INVX3 U240 ( .A(n235), .Y(n232) );
  INVX3 U241 ( .A(n234), .Y(n233) );
  CLKINVX1 U242 ( .A(n337), .Y(n250) );
  CLKINVX1 U243 ( .A(n352), .Y(n251) );
  CLKINVX1 U244 ( .A(n277), .Y(n252) );
  CLKBUFX3 U245 ( .A(SH[0]), .Y(n225) );
  CLKBUFX3 U246 ( .A(SH[0]), .Y(n226) );
  CLKBUFX3 U247 ( .A(n235), .Y(n234) );
  CLKBUFX3 U248 ( .A(SH[4]), .Y(n236) );
  CLKBUFX3 U249 ( .A(SH[4]), .Y(n237) );
  CLKINVX1 U250 ( .A(n288), .Y(n255) );
  CLKINVX1 U251 ( .A(n295), .Y(n242) );
  CLKBUFX3 U252 ( .A(SH[1]), .Y(n227) );
  CLKBUFX3 U253 ( .A(SH[2]), .Y(n230) );
  CLKINVX1 U254 ( .A(SH[3]), .Y(n235) );
  INVXL U255 ( .A(A[2]), .Y(n256) );
  CLKINVX1 U256 ( .A(n281), .Y(n254) );
  INVXL U257 ( .A(A[1]), .Y(n257) );
  MX3XL U258 ( .A(n261), .B(n262), .C(n240), .S0(n233), .S1(n237), .Y(B[8]) );
  MXI2X1 U259 ( .A(n264), .B(n265), .S0(n236), .Y(B[7]) );
  MX3XL U260 ( .A(n266), .B(n267), .C(n268), .S0(n230), .S1(n232), .Y(n264) );
  MXI2X1 U261 ( .A(n269), .B(n270), .S0(n236), .Y(B[6]) );
  MX3XL U262 ( .A(n271), .B(n272), .C(n273), .S0(n230), .S1(n232), .Y(n269) );
  MXI2X1 U263 ( .A(n274), .B(n275), .S0(n236), .Y(B[5]) );
  MX3XL U264 ( .A(n276), .B(n277), .C(n278), .S0(n230), .S1(n232), .Y(n274) );
  MXI2X1 U265 ( .A(n279), .B(n280), .S0(n236), .Y(B[4]) );
  MX3XL U266 ( .A(n281), .B(n282), .C(n283), .S0(n230), .S1(n232), .Y(n279) );
  MX3XL U267 ( .A(n287), .B(n288), .C(n266), .S0(n227), .S1(n230), .Y(n284) );
  MXI2X1 U268 ( .A(n289), .B(n290), .S0(n227), .Y(n266) );
  NOR2X1 U269 ( .A(SH[4]), .B(n291), .Y(B[31]) );
  NOR2X1 U270 ( .A(SH[4]), .B(n292), .Y(B[30]) );
  MX3XL U271 ( .A(n293), .B(n294), .C(n242), .S0(n233), .S1(n237), .Y(B[2]) );
  MX3XL U272 ( .A(n296), .B(n297), .C(n253), .S0(n227), .S1(n230), .Y(n293) );
  MXI2X1 U273 ( .A(n298), .B(n299), .S0(n227), .Y(n271) );
  NOR2X1 U274 ( .A(SH[4]), .B(n300), .Y(B[29]) );
  NOR2X1 U275 ( .A(n236), .B(n301), .Y(B[28]) );
  NOR2X1 U276 ( .A(n237), .B(n302), .Y(B[27]) );
  NOR2X1 U277 ( .A(n237), .B(n303), .Y(B[26]) );
  NOR2X1 U278 ( .A(n237), .B(n260), .Y(B[25]) );
  NAND2X1 U279 ( .A(n304), .B(n234), .Y(n260) );
  NOR2X1 U280 ( .A(n237), .B(n263), .Y(B[24]) );
  NOR2X1 U281 ( .A(n237), .B(n265), .Y(B[23]) );
  MXI2X1 U282 ( .A(n243), .B(n306), .S0(n232), .Y(n265) );
  MXI2X1 U283 ( .A(n244), .B(n308), .S0(n232), .Y(n270) );
  MXI2X1 U284 ( .A(n245), .B(n310), .S0(n232), .Y(n275) );
  NOR2X1 U285 ( .A(n237), .B(n280), .Y(B[20]) );
  MXI2X1 U286 ( .A(n246), .B(n312), .S0(n232), .Y(n280) );
  MXI2X1 U287 ( .A(n314), .B(n315), .S0(n236), .Y(B[1]) );
  MX3XL U288 ( .A(n316), .B(n276), .C(n258), .S0(n230), .S1(n232), .Y(n314) );
  MXI2X1 U289 ( .A(n252), .B(n317), .S0(n230), .Y(n258) );
  MXI2X1 U290 ( .A(n290), .B(n318), .S0(n227), .Y(n277) );
  MXI2X1 U291 ( .A(n255), .B(n289), .S0(n227), .Y(n276) );
  MX3XL U292 ( .A(n257), .B(n256), .C(n287), .S0(SH[0]), .S1(n227), .Y(n316)
         );
  NOR2X1 U293 ( .A(n237), .B(n285), .Y(B[19]) );
  MXI2X1 U294 ( .A(n319), .B(n320), .S0(n232), .Y(n285) );
  NOR2X1 U295 ( .A(n237), .B(n295), .Y(B[18]) );
  MXI2X1 U296 ( .A(n321), .B(n322), .S0(n232), .Y(n295) );
  NOR2X1 U297 ( .A(SH[4]), .B(n315), .Y(B[17]) );
  MXI2X1 U298 ( .A(n247), .B(n304), .S0(n232), .Y(n315) );
  MXI2X1 U299 ( .A(n325), .B(n326), .S0(n231), .Y(n259) );
  NOR2X1 U300 ( .A(n236), .B(n327), .Y(B[16]) );
  NOR2BX1 U301 ( .AN(n328), .B(n230), .Y(n306) );
  MXI2X1 U302 ( .A(n249), .B(n331), .S0(n230), .Y(n268) );
  NAND2X1 U303 ( .A(n308), .B(n234), .Y(n292) );
  NOR2BX1 U304 ( .AN(n333), .B(n230), .Y(n308) );
  MXI2X1 U305 ( .A(n334), .B(n335), .S0(n231), .Y(n309) );
  MXI2X1 U306 ( .A(n250), .B(n336), .S0(n230), .Y(n273) );
  NAND2X1 U307 ( .A(n310), .B(n234), .Y(n300) );
  CLKMX2X2 U308 ( .A(n338), .B(n339), .S0(n228), .Y(n323) );
  MXI2X1 U309 ( .A(n324), .B(n325), .S0(n231), .Y(n311) );
  CLKMX2X2 U310 ( .A(n340), .B(n341), .S0(n228), .Y(n325) );
  CLKMX2X2 U311 ( .A(n342), .B(n343), .S0(n229), .Y(n324) );
  MXI2X1 U312 ( .A(n317), .B(n326), .S0(n230), .Y(n278) );
  CLKMX2X2 U313 ( .A(n344), .B(n345), .S0(n229), .Y(n326) );
  CLKMX2X2 U314 ( .A(n346), .B(n347), .S0(n228), .Y(n317) );
  NAND2X1 U315 ( .A(n312), .B(n234), .Y(n301) );
  NOR2BX1 U316 ( .AN(n348), .B(n230), .Y(n312) );
  MXI2X1 U317 ( .A(n349), .B(n350), .S0(n231), .Y(n313) );
  MXI2X1 U318 ( .A(n251), .B(n351), .S0(n230), .Y(n283) );
  MX3XL U319 ( .A(n286), .B(n319), .C(n238), .S0(n233), .S1(n236), .Y(B[11])
         );
  CLKMX2X2 U320 ( .A(n328), .B(n329), .S0(n231), .Y(n320) );
  CLKMX2X2 U321 ( .A(n339), .B(n342), .S0(n228), .Y(n329) );
  NOR2BX1 U322 ( .AN(n338), .B(n227), .Y(n328) );
  CLKMX2X2 U323 ( .A(n330), .B(n331), .S0(n231), .Y(n319) );
  CLKMX2X2 U324 ( .A(n341), .B(n344), .S0(n228), .Y(n331) );
  CLKMX2X2 U325 ( .A(n343), .B(n340), .S0(n228), .Y(n330) );
  MXI2X1 U326 ( .A(n332), .B(n267), .S0(n231), .Y(n286) );
  MXI2X1 U327 ( .A(n318), .B(n347), .S0(n227), .Y(n267) );
  MXI2X1 U328 ( .A(n345), .B(n346), .S0(n229), .Y(n332) );
  MX3XL U329 ( .A(n294), .B(n321), .C(n241), .S0(n233), .S1(n236), .Y(B[10])
         );
  CLKMX2X2 U330 ( .A(n333), .B(n334), .S0(n231), .Y(n322) );
  CLKMX2X2 U331 ( .A(n353), .B(n354), .S0(n228), .Y(n334) );
  NOR2BX1 U332 ( .AN(n355), .B(n227), .Y(n333) );
  CLKMX2X2 U333 ( .A(n335), .B(n336), .S0(n231), .Y(n321) );
  CLKMX2X2 U334 ( .A(n356), .B(n357), .S0(n228), .Y(n336) );
  CLKMX2X2 U335 ( .A(n358), .B(n359), .S0(n228), .Y(n335) );
  MXI2X1 U336 ( .A(n337), .B(n272), .S0(n231), .Y(n294) );
  MXI2X1 U337 ( .A(n360), .B(n361), .S0(n227), .Y(n272) );
  MXI2X1 U338 ( .A(n362), .B(n363), .S0(n229), .Y(n337) );
  MX3XL U339 ( .A(n364), .B(n261), .C(n239), .S0(n233), .S1(n236), .Y(B[0]) );
  MXI2X1 U340 ( .A(n262), .B(n305), .S0(n232), .Y(n327) );
  CLKMX2X2 U341 ( .A(n348), .B(n349), .S0(n231), .Y(n305) );
  CLKMX2X2 U342 ( .A(n354), .B(n358), .S0(n228), .Y(n349) );
  CLKMX2X2 U343 ( .A(n355), .B(n353), .S0(n228), .Y(n348) );
  CLKMX2X2 U344 ( .A(n350), .B(n351), .S0(n231), .Y(n262) );
  CLKMX2X2 U345 ( .A(n357), .B(n362), .S0(n228), .Y(n351) );
  CLKMX2X2 U346 ( .A(n359), .B(n356), .S0(n228), .Y(n350) );
  MXI2X1 U347 ( .A(n352), .B(n282), .S0(n231), .Y(n261) );
  MXI2X1 U348 ( .A(n299), .B(n360), .S0(n227), .Y(n282) );
  MXI2X1 U349 ( .A(n363), .B(n361), .S0(n229), .Y(n352) );
  MX3XL U350 ( .A(n365), .B(n296), .C(n254), .S0(n227), .S1(n230), .Y(n364) );
  MXI2X1 U351 ( .A(n297), .B(n298), .S0(n227), .Y(n281) );
endmodule


module Execution_DW_leftsh_0 ( A, SH, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  wire   n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360;

  MXI3X1 U178 ( .A(n291), .B(n326), .C(n272), .S0(n231), .S1(n234), .Y(B[18])
         );
  MXI3X1 U179 ( .A(n303), .B(n301), .C(n335), .S0(n231), .S1(n234), .Y(B[16])
         );
  MXI3X1 U180 ( .A(n297), .B(n295), .C(n321), .S0(n231), .S1(n235), .Y(B[17])
         );
  MXI3X1 U181 ( .A(n286), .B(n322), .C(n260), .S0(n231), .S1(n235), .Y(B[19])
         );
  MXI3X1 U182 ( .A(n270), .B(n309), .C(n257), .S0(n231), .S1(n234), .Y(B[22])
         );
  MXI3X1 U183 ( .A(A[30]), .B(A[29]), .C(n271), .S0(SH[0]), .S1(SH[1]), .Y(
        n222) );
  MX2X1 U184 ( .A(n344), .B(n345), .S0(n229), .Y(n310) );
  CLKMX2X2 U185 ( .A(n354), .B(n336), .S0(n229), .Y(n318) );
  NOR2BX1 U186 ( .AN(n354), .B(n228), .Y(n300) );
  MX2X1 U187 ( .A(n340), .B(n341), .S0(n229), .Y(n306) );
  INVX1 U188 ( .A(n309), .Y(n244) );
  MX2XL U189 ( .A(A[14]), .B(A[13]), .S0(n224), .Y(n339) );
  NOR2BX1 U190 ( .AN(n344), .B(SH[2]), .Y(n327) );
  NOR2BX1 U191 ( .AN(n340), .B(n228), .Y(n323) );
  MX2XL U192 ( .A(A[1]), .B(A[0]), .S0(n223), .Y(n350) );
  MXI2XL U193 ( .A(n319), .B(n302), .S0(n229), .Y(n279) );
  MXI2XL U194 ( .A(n315), .B(n296), .S0(n229), .Y(n274) );
  MX2X1 U195 ( .A(n330), .B(n331), .S0(n229), .Y(n314) );
  NOR2X1 U196 ( .A(n235), .B(n284), .Y(B[11]) );
  NOR2X1 U197 ( .A(n235), .B(n289), .Y(B[10]) );
  NOR2X1 U198 ( .A(SH[4]), .B(n255), .Y(B[8]) );
  NOR2BX1 U199 ( .AN(n330), .B(n228), .Y(n294) );
  NOR2XL U200 ( .A(n235), .B(n268), .Y(B[14]) );
  NOR2XL U201 ( .A(n235), .B(n263), .Y(B[15]) );
  NOR2XL U202 ( .A(n235), .B(n280), .Y(B[12]) );
  NOR2XL U203 ( .A(n235), .B(n272), .Y(B[2]) );
  NOR2XL U204 ( .A(n235), .B(n335), .Y(B[0]) );
  NOR2XL U205 ( .A(n235), .B(n275), .Y(B[13]) );
  NOR2XL U206 ( .A(n235), .B(n254), .Y(B[9]) );
  NOR2XL U207 ( .A(n235), .B(n321), .Y(B[1]) );
  NOR2XL U208 ( .A(n235), .B(n260), .Y(B[3]) );
  NOR2XL U209 ( .A(n235), .B(n259), .Y(B[4]) );
  NOR2XL U210 ( .A(n235), .B(n256), .Y(B[7]) );
  NOR2XL U211 ( .A(n235), .B(n257), .Y(B[6]) );
  NOR2XL U212 ( .A(n235), .B(n258), .Y(B[5]) );
  NOR2BXL U213 ( .AN(A[0]), .B(SH[0]), .Y(n360) );
  MX2XL U214 ( .A(A[9]), .B(A[8]), .S0(n224), .Y(n353) );
  MX2XL U215 ( .A(A[13]), .B(A[12]), .S0(n223), .Y(n343) );
  MX2XL U216 ( .A(A[11]), .B(A[10]), .S0(n223), .Y(n351) );
  MX2XL U217 ( .A(A[8]), .B(A[7]), .S0(n223), .Y(n359) );
  MX2XL U218 ( .A(A[10]), .B(A[9]), .S0(n223), .Y(n357) );
  MX2XL U219 ( .A(A[12]), .B(A[11]), .S0(n223), .Y(n347) );
  MX2XL U220 ( .A(A[3]), .B(A[2]), .S0(n223), .Y(n348) );
  MX2XL U221 ( .A(A[4]), .B(A[3]), .S0(n223), .Y(n356) );
  MX2XL U222 ( .A(A[6]), .B(A[5]), .S0(n223), .Y(n358) );
  MX2XL U223 ( .A(A[7]), .B(A[6]), .S0(n223), .Y(n352) );
  MX2XL U224 ( .A(A[2]), .B(A[1]), .S0(n223), .Y(n355) );
  MX2XL U225 ( .A(A[5]), .B(A[4]), .S0(n223), .Y(n349) );
  MX2XL U226 ( .A(A[16]), .B(A[15]), .S0(n224), .Y(n329) );
  MX2XL U227 ( .A(A[15]), .B(A[14]), .S0(n224), .Y(n334) );
  MX2XL U228 ( .A(A[18]), .B(A[17]), .S0(n224), .Y(n320) );
  MX2XL U229 ( .A(A[17]), .B(A[16]), .S0(n224), .Y(n325) );
  MX2XL U230 ( .A(A[19]), .B(A[18]), .S0(n224), .Y(n316) );
  MX2XL U231 ( .A(A[22]), .B(A[21]), .S0(n224), .Y(n304) );
  MX2XL U232 ( .A(A[20]), .B(A[19]), .S0(n224), .Y(n312) );
  MX2XL U233 ( .A(A[25]), .B(A[24]), .S0(n224), .Y(n287) );
  MX2XL U234 ( .A(A[23]), .B(A[22]), .S0(n224), .Y(n298) );
  MX2XL U235 ( .A(A[21]), .B(A[20]), .S0(n224), .Y(n308) );
  MX2XL U236 ( .A(A[24]), .B(A[23]), .S0(n224), .Y(n292) );
  MX2XL U237 ( .A(A[27]), .B(A[26]), .S0(n224), .Y(n276) );
  MX2XL U238 ( .A(A[26]), .B(A[25]), .S0(n224), .Y(n281) );
  MX2XL U239 ( .A(A[28]), .B(A[27]), .S0(SH[0]), .Y(n271) );
  MX2XL U240 ( .A(A[29]), .B(A[28]), .S0(n224), .Y(n265) );
  MX2XL U241 ( .A(A[31]), .B(A[30]), .S0(n223), .Y(n264) );
  CLKINVX1 U242 ( .A(n263), .Y(n243) );
  CLKINVX1 U243 ( .A(n280), .Y(n246) );
  CLKINVX1 U244 ( .A(n275), .Y(n245) );
  CLKINVX1 U245 ( .A(n322), .Y(n247) );
  CLKINVX1 U246 ( .A(n326), .Y(n248) );
  CLKINVX1 U247 ( .A(n295), .Y(n249) );
  CLKINVX1 U248 ( .A(n301), .Y(n250) );
  INVX3 U249 ( .A(n225), .Y(n226) );
  INVX3 U250 ( .A(n228), .Y(n229) );
  INVX3 U251 ( .A(n233), .Y(n230) );
  INVX3 U252 ( .A(n232), .Y(n231) );
  CLKINVX1 U253 ( .A(n225), .Y(n227) );
  CLKINVX1 U254 ( .A(n307), .Y(n240) );
  CLKINVX1 U255 ( .A(n315), .Y(n241) );
  CLKINVX1 U256 ( .A(n319), .Y(n242) );
  CLKINVX1 U257 ( .A(n290), .Y(n239) );
  CLKINVX1 U258 ( .A(n266), .Y(n236) );
  CLKINVX1 U259 ( .A(n277), .Y(n237) );
  CLKINVX1 U260 ( .A(n258), .Y(n252) );
  CLKINVX1 U261 ( .A(n256), .Y(n251) );
  CLKINVX1 U262 ( .A(n259), .Y(n253) );
  CLKBUFX3 U263 ( .A(SH[0]), .Y(n223) );
  CLKBUFX3 U264 ( .A(SH[0]), .Y(n224) );
  CLKBUFX3 U265 ( .A(n233), .Y(n232) );
  CLKBUFX3 U266 ( .A(SH[4]), .Y(n234) );
  CLKBUFX3 U267 ( .A(SH[4]), .Y(n235) );
  CLKINVX1 U268 ( .A(n282), .Y(n238) );
  CLKBUFX3 U269 ( .A(SH[2]), .Y(n228) );
  CLKBUFX3 U270 ( .A(SH[1]), .Y(n225) );
  CLKINVX1 U271 ( .A(SH[3]), .Y(n233) );
  MX3XL U272 ( .A(n261), .B(n262), .C(n243), .S0(n231), .S1(n234), .Y(B[31])
         );
  MX3XL U273 ( .A(n264), .B(n265), .C(n236), .S0(n225), .S1(n228), .Y(n261) );
  MXI2X1 U274 ( .A(n267), .B(n268), .S0(n234), .Y(B[30]) );
  MX3XL U275 ( .A(n222), .B(n269), .C(n270), .S0(n228), .S1(n230), .Y(n267) );
  MX3XL U276 ( .A(n273), .B(n274), .C(n245), .S0(n231), .S1(n234), .Y(B[29])
         );
  MX3XL U277 ( .A(n265), .B(n276), .C(n237), .S0(n225), .S1(n228), .Y(n273) );
  MX3XL U278 ( .A(n278), .B(n279), .C(n246), .S0(n231), .S1(n234), .Y(B[28])
         );
  MX3XL U279 ( .A(n271), .B(n281), .C(n238), .S0(n225), .S1(n228), .Y(n278) );
  MXI2X1 U280 ( .A(n283), .B(n284), .S0(n234), .Y(B[27]) );
  MX3XL U281 ( .A(n266), .B(n285), .C(n286), .S0(n228), .S1(n230), .Y(n283) );
  MXI2X1 U282 ( .A(n276), .B(n287), .S0(n225), .Y(n266) );
  MXI2X1 U283 ( .A(n288), .B(n289), .S0(n234), .Y(B[26]) );
  MX3XL U284 ( .A(n269), .B(n290), .C(n291), .S0(n228), .S1(n230), .Y(n288) );
  MXI2X1 U285 ( .A(n281), .B(n292), .S0(n225), .Y(n269) );
  MXI2X1 U286 ( .A(n293), .B(n254), .S0(n234), .Y(B[25]) );
  MXI2X1 U287 ( .A(n249), .B(n294), .S0(n230), .Y(n254) );
  MX3XL U288 ( .A(n277), .B(n296), .C(n297), .S0(n228), .S1(n230), .Y(n293) );
  MXI2X1 U289 ( .A(n287), .B(n298), .S0(n225), .Y(n277) );
  MXI2X1 U290 ( .A(n299), .B(n255), .S0(n234), .Y(B[24]) );
  MXI2X1 U291 ( .A(n250), .B(n300), .S0(n230), .Y(n255) );
  MX3XL U292 ( .A(n282), .B(n302), .C(n303), .S0(n228), .S1(n230), .Y(n299) );
  MXI2X1 U293 ( .A(n292), .B(n304), .S0(n225), .Y(n282) );
  MX3XL U294 ( .A(n262), .B(n305), .C(n251), .S0(n231), .S1(n234), .Y(B[23])
         );
  NAND2X1 U295 ( .A(n306), .B(n232), .Y(n256) );
  MXI2X1 U296 ( .A(n307), .B(n285), .S0(n229), .Y(n262) );
  MXI2X1 U297 ( .A(n298), .B(n308), .S0(n225), .Y(n285) );
  NAND2X1 U298 ( .A(n310), .B(n232), .Y(n257) );
  MXI2X1 U299 ( .A(n239), .B(n311), .S0(n228), .Y(n270) );
  MXI2X1 U300 ( .A(n304), .B(n312), .S0(n225), .Y(n290) );
  MX3XL U301 ( .A(n274), .B(n313), .C(n252), .S0(n231), .S1(n234), .Y(B[21])
         );
  NAND2X1 U302 ( .A(n314), .B(n232), .Y(n258) );
  MXI2X1 U303 ( .A(n308), .B(n316), .S0(n225), .Y(n296) );
  MX3XL U304 ( .A(n279), .B(n317), .C(n253), .S0(n231), .S1(n235), .Y(B[20])
         );
  NAND2X1 U305 ( .A(n318), .B(n232), .Y(n259) );
  MXI2X1 U306 ( .A(n312), .B(n320), .S0(n225), .Y(n302) );
  NAND2X1 U307 ( .A(n323), .B(n232), .Y(n260) );
  MXI2X1 U308 ( .A(n240), .B(n324), .S0(n228), .Y(n286) );
  MXI2X1 U309 ( .A(n325), .B(n316), .S0(n227), .Y(n307) );
  NAND2X1 U310 ( .A(n327), .B(n232), .Y(n272) );
  MXI2X1 U311 ( .A(n311), .B(n328), .S0(n228), .Y(n291) );
  CLKMX2X2 U312 ( .A(n329), .B(n320), .S0(n227), .Y(n311) );
  NAND2X1 U313 ( .A(n294), .B(n232), .Y(n321) );
  MXI2X1 U314 ( .A(n331), .B(n332), .S0(n229), .Y(n295) );
  MXI2X1 U315 ( .A(n241), .B(n333), .S0(n228), .Y(n297) );
  MXI2X1 U316 ( .A(n334), .B(n325), .S0(n227), .Y(n315) );
  MXI2X1 U317 ( .A(n336), .B(n337), .S0(n229), .Y(n301) );
  MXI2X1 U318 ( .A(n242), .B(n338), .S0(n228), .Y(n303) );
  MXI2X1 U319 ( .A(n339), .B(n329), .S0(n227), .Y(n319) );
  MXI2X1 U320 ( .A(n305), .B(n306), .S0(n230), .Y(n263) );
  CLKMX2X2 U321 ( .A(n342), .B(n324), .S0(n229), .Y(n305) );
  CLKMX2X2 U322 ( .A(n343), .B(n334), .S0(n227), .Y(n324) );
  MXI2X1 U323 ( .A(n244), .B(n310), .S0(n230), .Y(n268) );
  MXI2X1 U324 ( .A(n346), .B(n328), .S0(n229), .Y(n309) );
  CLKMX2X2 U325 ( .A(n347), .B(n339), .S0(n226), .Y(n328) );
  MXI2X1 U326 ( .A(n313), .B(n314), .S0(n230), .Y(n275) );
  CLKMX2X2 U327 ( .A(n348), .B(n349), .S0(n226), .Y(n331) );
  NOR2BX1 U328 ( .AN(n350), .B(n225), .Y(n330) );
  CLKMX2X2 U329 ( .A(n332), .B(n333), .S0(n229), .Y(n313) );
  CLKMX2X2 U330 ( .A(n351), .B(n343), .S0(n226), .Y(n333) );
  CLKMX2X2 U331 ( .A(n352), .B(n353), .S0(n226), .Y(n332) );
  MXI2X1 U332 ( .A(n317), .B(n318), .S0(n230), .Y(n280) );
  CLKMX2X2 U333 ( .A(n355), .B(n356), .S0(n226), .Y(n336) );
  CLKMX2X2 U334 ( .A(n337), .B(n338), .S0(n229), .Y(n317) );
  CLKMX2X2 U335 ( .A(n357), .B(n347), .S0(n226), .Y(n338) );
  CLKMX2X2 U336 ( .A(n358), .B(n359), .S0(n226), .Y(n337) );
  MXI2X1 U337 ( .A(n247), .B(n323), .S0(n230), .Y(n284) );
  CLKMX2X2 U338 ( .A(n350), .B(n348), .S0(n226), .Y(n340) );
  MXI2X1 U339 ( .A(n341), .B(n342), .S0(n229), .Y(n322) );
  CLKMX2X2 U340 ( .A(n353), .B(n351), .S0(n226), .Y(n342) );
  CLKMX2X2 U341 ( .A(n349), .B(n352), .S0(n226), .Y(n341) );
  MXI2X1 U342 ( .A(n248), .B(n327), .S0(n230), .Y(n289) );
  CLKMX2X2 U343 ( .A(n360), .B(n355), .S0(n226), .Y(n344) );
  MXI2X1 U344 ( .A(n345), .B(n346), .S0(n229), .Y(n326) );
  CLKMX2X2 U345 ( .A(n359), .B(n357), .S0(n226), .Y(n346) );
  CLKMX2X2 U346 ( .A(n356), .B(n358), .S0(n226), .Y(n345) );
  NAND2X1 U347 ( .A(n300), .B(n232), .Y(n335) );
  NOR2BX1 U348 ( .AN(n360), .B(n225), .Y(n354) );
endmodule


module Execution_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n34, n36, n38, n39, n40, n41, n42, n44, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n60, n62, n63, n64, n65,
         n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n127, n128, n129, n130,
         n132, n133, n134, n135, n136, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374;

  OAI21X2 U298 ( .A0(n66), .A1(n70), .B0(n67), .Y(n65) );
  OAI21XL U299 ( .A0(n171), .A1(n175), .B0(n172), .Y(n170) );
  CLKINVX1 U300 ( .A(B[20]), .Y(n242) );
  CLKINVX1 U301 ( .A(B[21]), .Y(n241) );
  NOR2X1 U302 ( .A(n174), .B(n171), .Y(n169) );
  CLKINVX1 U303 ( .A(B[17]), .Y(n245) );
  CLKINVX1 U304 ( .A(B[19]), .Y(n243) );
  CLKINVX1 U305 ( .A(B[23]), .Y(n239) );
  CLKINVX1 U306 ( .A(B[25]), .Y(n237) );
  CLKINVX1 U307 ( .A(B[24]), .Y(n238) );
  CLKINVX1 U308 ( .A(B[22]), .Y(n240) );
  OAI21XL U309 ( .A0(n87), .A1(n91), .B0(n88), .Y(n86) );
  OAI21XL U310 ( .A0(n197), .A1(n199), .B0(n198), .Y(n196) );
  OAI21XL U311 ( .A0(n179), .A1(n185), .B0(n180), .Y(n178) );
  CLKINVX1 U312 ( .A(B[13]), .Y(n249) );
  OAI21XL U313 ( .A0(n135), .A1(n141), .B0(n136), .Y(n134) );
  NOR2X1 U314 ( .A(n57), .B(n52), .Y(n50) );
  NOR2X1 U315 ( .A(n253), .B(A[9]), .Y(n160) );
  NOR2X1 U316 ( .A(n247), .B(A[15]), .Y(n123) );
  NAND2X1 U317 ( .A(n260), .B(A[2]), .Y(n194) );
  NOR2X1 U318 ( .A(n251), .B(A[11]), .Y(n148) );
  NOR2X1 U319 ( .A(n140), .B(n135), .Y(n133) );
  INVX1 U320 ( .A(B[7]), .Y(n255) );
  INVX1 U321 ( .A(B[2]), .Y(n260) );
  NOR2X1 U322 ( .A(n144), .B(n119), .Y(n117) );
  AOI21X2 U323 ( .A0(n159), .A1(n146), .B0(n147), .Y(n145) );
  NOR2X1 U324 ( .A(n237), .B(A[25]), .Y(n66) );
  NOR2X1 U325 ( .A(n243), .B(A[19]), .Y(n100) );
  INVXL U326 ( .A(B[0]), .Y(n262) );
  NOR2X1 U327 ( .A(n241), .B(A[21]), .Y(n87) );
  NAND2XL U328 ( .A(n247), .B(A[15]), .Y(n124) );
  INVXL U329 ( .A(B[16]), .Y(n246) );
  INVXL U330 ( .A(B[27]), .Y(n235) );
  INVX1 U331 ( .A(B[26]), .Y(n236) );
  INVX1 U332 ( .A(B[18]), .Y(n244) );
  CLKINVX4 U333 ( .A(n142), .Y(n365) );
  NAND2X4 U334 ( .A(n366), .B(n132), .Y(n130) );
  AOI21X2 U335 ( .A0(n166), .A1(n117), .B0(n118), .Y(n116) );
  OAI21X1 U336 ( .A0(n116), .A1(n48), .B0(n49), .Y(n47) );
  XNOR2X1 U337 ( .A(n130), .B(n18), .Y(DIFF[14]) );
  AO21X2 U338 ( .A0(n130), .A1(n217), .B0(n127), .Y(n368) );
  XNOR2X4 U339 ( .A(n368), .B(n17), .Y(DIFF[15]) );
  NAND2X1 U340 ( .A(n252), .B(A[10]), .Y(n154) );
  INVX1 U341 ( .A(n143), .Y(n142) );
  NAND2X1 U342 ( .A(n365), .B(n133), .Y(n366) );
  CLKINVX1 U343 ( .A(B[1]), .Y(n261) );
  INVXL U344 ( .A(n134), .Y(n132) );
  NAND2XL U345 ( .A(n255), .B(A[7]), .Y(n172) );
  AOI21XL U346 ( .A0(n115), .A1(n106), .B0(n107), .Y(n105) );
  INVX1 U347 ( .A(n159), .Y(n157) );
  INVXL U348 ( .A(n158), .Y(n156) );
  NOR2X1 U349 ( .A(n255), .B(A[7]), .Y(n171) );
  AOI21X2 U350 ( .A0(n115), .A1(n94), .B0(n95), .Y(n93) );
  NOR2X1 U351 ( .A(n163), .B(n160), .Y(n158) );
  OR2X1 U352 ( .A(n160), .B(n164), .Y(n367) );
  NAND2X1 U353 ( .A(n367), .B(n161), .Y(n159) );
  NAND2X1 U354 ( .A(n258), .B(A[4]), .Y(n185) );
  NOR2X1 U355 ( .A(n260), .B(A[2]), .Y(n193) );
  NAND2XL U356 ( .A(n245), .B(A[17]), .Y(n109) );
  NOR2X1 U357 ( .A(n239), .B(A[23]), .Y(n79) );
  NOR2X1 U358 ( .A(n240), .B(A[22]), .Y(n82) );
  NAND2XL U359 ( .A(n251), .B(A[11]), .Y(n149) );
  NAND2XL U360 ( .A(n242), .B(A[20]), .Y(n91) );
  NAND2XL U361 ( .A(n240), .B(A[22]), .Y(n83) );
  NAND2X1 U362 ( .A(n238), .B(A[24]), .Y(n70) );
  NOR2XL U363 ( .A(n233), .B(A[29]), .Y(n40) );
  NAND2XL U364 ( .A(n254), .B(A[8]), .Y(n164) );
  CLKINVX1 U365 ( .A(B[8]), .Y(n254) );
  NAND2XL U366 ( .A(n253), .B(A[9]), .Y(n161) );
  OAI21XL U367 ( .A0(n165), .A1(n144), .B0(n145), .Y(n143) );
  AOI21X1 U368 ( .A0(n92), .A1(n85), .B0(n86), .Y(n84) );
  AOI21X1 U369 ( .A0(n115), .A1(n73), .B0(n74), .Y(n72) );
  INVXL U370 ( .A(n97), .Y(n95) );
  INVXL U371 ( .A(n187), .Y(n186) );
  AO21X1 U372 ( .A0(n155), .A1(n221), .B0(n152), .Y(n370) );
  OAI21X1 U373 ( .A0(n108), .A1(n114), .B0(n109), .Y(n107) );
  NAND2XL U374 ( .A(n373), .B(n46), .Y(n4) );
  NAND2X1 U375 ( .A(n64), .B(n371), .Y(n57) );
  XOR2X1 U376 ( .A(n176), .B(n26), .Y(DIFF[6]) );
  INVXL U377 ( .A(n163), .Y(n223) );
  NAND2X1 U378 ( .A(n261), .B(A[1]), .Y(n198) );
  NOR2X1 U379 ( .A(n249), .B(A[13]), .Y(n135) );
  INVXL U380 ( .A(B[28]), .Y(n234) );
  NOR2X2 U381 ( .A(n75), .B(n96), .Y(n73) );
  OAI21X1 U382 ( .A0(n145), .A1(n119), .B0(n120), .Y(n118) );
  NAND2X2 U383 ( .A(n133), .B(n121), .Y(n119) );
  INVXL U384 ( .A(n96), .Y(n94) );
  NAND2XL U385 ( .A(n158), .B(n146), .Y(n144) );
  INVXL U386 ( .A(n58), .Y(n56) );
  XNOR2XL U387 ( .A(n92), .B(n12), .Y(DIFF[20]) );
  XOR2XL U388 ( .A(n84), .B(n10), .Y(DIFF[22]) );
  XNOR2XL U389 ( .A(n71), .B(n8), .Y(DIFF[24]) );
  AOI21XL U390 ( .A0(n186), .A1(n177), .B0(n178), .Y(n176) );
  XOR2XL U391 ( .A(n105), .B(n14), .Y(DIFF[18]) );
  OAI21X1 U392 ( .A0(n42), .A1(n40), .B0(n41), .Y(n39) );
  OAI21X2 U393 ( .A0(n97), .A1(n75), .B0(n76), .Y(n74) );
  OAI21X2 U394 ( .A0(n187), .A1(n167), .B0(n168), .Y(n166) );
  NAND2XL U395 ( .A(n217), .B(n129), .Y(n18) );
  XNOR2XL U396 ( .A(n39), .B(n2), .Y(DIFF[30]) );
  INVXL U397 ( .A(n160), .Y(n222) );
  NAND2XL U398 ( .A(n225), .B(n175), .Y(n26) );
  INVXL U399 ( .A(n174), .Y(n225) );
  XOR2XL U400 ( .A(n142), .B(n20), .Y(DIFF[12]) );
  NAND2XL U401 ( .A(n219), .B(n141), .Y(n20) );
  XOR2XL U402 ( .A(n165), .B(n24), .Y(DIFF[8]) );
  XNOR2X1 U403 ( .A(n369), .B(n19), .Y(DIFF[13]) );
  AO21XL U404 ( .A0(n143), .A1(n219), .B0(n139), .Y(n369) );
  XNOR2X1 U405 ( .A(n370), .B(n21), .Y(DIFF[11]) );
  AOI21XL U406 ( .A0(n115), .A1(n215), .B0(n112), .Y(n110) );
  INVXL U407 ( .A(n114), .Y(n112) );
  NAND2XL U408 ( .A(n215), .B(n114), .Y(n16) );
  XNOR2XL U409 ( .A(n115), .B(n16), .Y(DIFF[16]) );
  XNOR2XL U410 ( .A(n47), .B(n4), .Y(DIFF[28]) );
  XOR2XL U411 ( .A(n42), .B(n3), .Y(DIFF[29]) );
  XOR2XL U412 ( .A(n31), .B(n199), .Y(DIFF[1]) );
  INVXL U413 ( .A(n197), .Y(n230) );
  XOR2XL U414 ( .A(n195), .B(n30), .Y(DIFF[2]) );
  AOI21XL U415 ( .A0(n186), .A1(n227), .B0(n183), .Y(n181) );
  INVXL U416 ( .A(n179), .Y(n226) );
  XNOR2XL U417 ( .A(n186), .B(n28), .Y(DIFF[4]) );
  NAND2XL U418 ( .A(n227), .B(n185), .Y(n28) );
  INVXL U419 ( .A(n190), .Y(n228) );
  INVXL U420 ( .A(n140), .Y(n219) );
  INVXL U421 ( .A(n153), .Y(n221) );
  INVXL U422 ( .A(n128), .Y(n217) );
  NAND2BXL U423 ( .AN(n69), .B(n70), .Y(n8) );
  NAND2BXL U424 ( .AN(n103), .B(n104), .Y(n14) );
  NAND2XL U425 ( .A(n371), .B(n62), .Y(n6) );
  INVXL U426 ( .A(n141), .Y(n139) );
  INVXL U427 ( .A(n129), .Y(n127) );
  NAND2XL U428 ( .A(n249), .B(A[13]), .Y(n136) );
  NAND2XL U429 ( .A(n259), .B(A[3]), .Y(n191) );
  NOR2XL U430 ( .A(n258), .B(A[4]), .Y(n184) );
  NOR2XL U431 ( .A(n246), .B(A[16]), .Y(n113) );
  NOR2X1 U432 ( .A(n245), .B(A[17]), .Y(n108) );
  NOR2X1 U433 ( .A(n254), .B(A[8]), .Y(n163) );
  NAND2XL U434 ( .A(n237), .B(A[25]), .Y(n67) );
  NAND2XL U435 ( .A(n241), .B(A[21]), .Y(n88) );
  NAND2XL U436 ( .A(n236), .B(A[26]), .Y(n62) );
  NAND2XL U437 ( .A(n257), .B(A[5]), .Y(n180) );
  NAND2XL U438 ( .A(n239), .B(A[23]), .Y(n80) );
  NAND2XL U439 ( .A(n235), .B(A[27]), .Y(n53) );
  NAND2XL U440 ( .A(n243), .B(A[19]), .Y(n101) );
  NOR2X1 U441 ( .A(n242), .B(A[20]), .Y(n90) );
  NOR2X1 U442 ( .A(n244), .B(A[18]), .Y(n103) );
  NOR2X1 U443 ( .A(n235), .B(A[27]), .Y(n52) );
  NAND2XL U444 ( .A(n232), .B(A[30]), .Y(n38) );
  NAND2XL U445 ( .A(n234), .B(A[28]), .Y(n46) );
  NAND2XL U446 ( .A(n233), .B(A[29]), .Y(n41) );
  OR2XL U447 ( .A(n232), .B(A[30]), .Y(n372) );
  OR2XL U448 ( .A(n234), .B(A[28]), .Y(n373) );
  INVXL U449 ( .A(B[29]), .Y(n233) );
  INVXL U450 ( .A(B[30]), .Y(n232) );
  INVXL U451 ( .A(B[31]), .Y(n231) );
  NOR2XL U452 ( .A(n231), .B(A[31]), .Y(n32) );
  AND2XL U453 ( .A(n231), .B(A[31]), .Y(n374) );
  XNOR2XL U454 ( .A(n262), .B(A[0]), .Y(DIFF[0]) );
  CLKINVX1 U455 ( .A(n116), .Y(n115) );
  CLKINVX1 U456 ( .A(n72), .Y(n71) );
  CLKINVX1 U457 ( .A(n93), .Y(n92) );
  OAI21XL U458 ( .A0(n165), .A1(n156), .B0(n157), .Y(n155) );
  CLKINVX1 U459 ( .A(n166), .Y(n165) );
  AOI21X1 U460 ( .A0(n71), .A1(n64), .B0(n65), .Y(n63) );
  AOI21X1 U461 ( .A0(n71), .A1(n55), .B0(n56), .Y(n54) );
  CLKINVX1 U462 ( .A(n57), .Y(n55) );
  NAND2X1 U463 ( .A(n77), .B(n85), .Y(n75) );
  XNOR2X1 U464 ( .A(n68), .B(n7), .Y(DIFF[25]) );
  XOR2X1 U465 ( .A(n63), .B(n6), .Y(DIFF[26]) );
  XOR2X1 U466 ( .A(n54), .B(n5), .Y(DIFF[27]) );
  XNOR2X1 U467 ( .A(n89), .B(n11), .Y(DIFF[21]) );
  XNOR2X1 U468 ( .A(n81), .B(n9), .Y(DIFF[23]) );
  XNOR2X1 U469 ( .A(n102), .B(n13), .Y(DIFF[19]) );
  CLKINVX1 U470 ( .A(n196), .Y(n195) );
  NAND2X1 U471 ( .A(n98), .B(n106), .Y(n96) );
  AOI21X1 U472 ( .A0(n47), .A1(n373), .B0(n44), .Y(n42) );
  CLKINVX1 U473 ( .A(n46), .Y(n44) );
  NAND2X1 U474 ( .A(n169), .B(n177), .Y(n167) );
  AOI21X1 U475 ( .A0(n178), .A1(n169), .B0(n170), .Y(n168) );
  AOI21X1 U476 ( .A0(n65), .A1(n371), .B0(n60), .Y(n58) );
  CLKINVX1 U477 ( .A(n62), .Y(n60) );
  AOI21X1 U478 ( .A0(n107), .A1(n98), .B0(n99), .Y(n97) );
  OAI21XL U479 ( .A0(n100), .A1(n104), .B0(n101), .Y(n99) );
  AOI21X1 U480 ( .A0(n196), .A1(n188), .B0(n189), .Y(n187) );
  OAI21XL U481 ( .A0(n190), .A1(n194), .B0(n191), .Y(n189) );
  NOR2X1 U482 ( .A(n193), .B(n190), .Y(n188) );
  AOI21X1 U483 ( .A0(n86), .A1(n77), .B0(n78), .Y(n76) );
  OAI21XL U484 ( .A0(n79), .A1(n83), .B0(n80), .Y(n78) );
  OAI21XL U485 ( .A0(n148), .A1(n154), .B0(n149), .Y(n147) );
  NAND2X1 U486 ( .A(n50), .B(n73), .Y(n48) );
  AOI21X1 U487 ( .A0(n74), .A1(n50), .B0(n51), .Y(n49) );
  XNOR2X1 U488 ( .A(n155), .B(n22), .Y(DIFF[10]) );
  NAND2X1 U489 ( .A(n221), .B(n154), .Y(n22) );
  XNOR2X1 U490 ( .A(n162), .B(n23), .Y(DIFF[9]) );
  NAND2X1 U491 ( .A(n222), .B(n161), .Y(n23) );
  OAI21XL U492 ( .A0(n165), .A1(n163), .B0(n164), .Y(n162) );
  XNOR2X1 U493 ( .A(n173), .B(n25), .Y(DIFF[7]) );
  NAND2X1 U494 ( .A(n224), .B(n172), .Y(n25) );
  OAI21XL U495 ( .A0(n176), .A1(n174), .B0(n175), .Y(n173) );
  CLKINVX1 U496 ( .A(n171), .Y(n224) );
  OAI21XL U497 ( .A0(n58), .A1(n52), .B0(n53), .Y(n51) );
  NOR2X1 U498 ( .A(n79), .B(n82), .Y(n77) );
  NOR2X1 U499 ( .A(n100), .B(n103), .Y(n98) );
  NOR2X1 U500 ( .A(n87), .B(n90), .Y(n85) );
  NOR2X1 U501 ( .A(n179), .B(n184), .Y(n177) );
  NOR2X1 U502 ( .A(n153), .B(n148), .Y(n146) );
  NOR2X1 U503 ( .A(n128), .B(n123), .Y(n121) );
  OAI21XL U504 ( .A0(n72), .A1(n69), .B0(n70), .Y(n68) );
  OAI21XL U505 ( .A0(n93), .A1(n90), .B0(n91), .Y(n89) );
  OAI21XL U506 ( .A0(n105), .A1(n103), .B0(n104), .Y(n102) );
  OAI21XL U507 ( .A0(n84), .A1(n82), .B0(n83), .Y(n81) );
  AOI21X1 U508 ( .A0(n39), .A1(n372), .B0(n36), .Y(n34) );
  CLKINVX1 U509 ( .A(n38), .Y(n36) );
  AOI21X1 U510 ( .A0(n134), .A1(n121), .B0(n122), .Y(n120) );
  OAI21XL U511 ( .A0(n123), .A1(n129), .B0(n124), .Y(n122) );
  XOR2X1 U512 ( .A(n34), .B(n1), .Y(DIFF[31]) );
  XOR2X1 U513 ( .A(n110), .B(n15), .Y(DIFF[17]) );
  NAND2X1 U514 ( .A(n214), .B(n109), .Y(n15) );
  XOR2X1 U515 ( .A(n181), .B(n27), .Y(DIFF[5]) );
  NAND2X1 U516 ( .A(n226), .B(n180), .Y(n27) );
  NAND2X1 U517 ( .A(n216), .B(n124), .Y(n17) );
  CLKINVX1 U518 ( .A(n123), .Y(n216) );
  NAND2X1 U519 ( .A(n220), .B(n149), .Y(n21) );
  CLKINVX1 U520 ( .A(n148), .Y(n220) );
  NAND2X1 U521 ( .A(n218), .B(n136), .Y(n19) );
  CLKINVX1 U522 ( .A(n135), .Y(n218) );
  NAND2X1 U523 ( .A(n223), .B(n164), .Y(n24) );
  XNOR2X1 U524 ( .A(n192), .B(n29), .Y(DIFF[3]) );
  NAND2X1 U525 ( .A(n228), .B(n191), .Y(n29) );
  OAI21XL U526 ( .A0(n195), .A1(n193), .B0(n194), .Y(n192) );
  NOR2X1 U527 ( .A(n108), .B(n113), .Y(n106) );
  NOR2X1 U528 ( .A(n69), .B(n66), .Y(n64) );
  CLKINVX1 U529 ( .A(n184), .Y(n227) );
  CLKINVX1 U530 ( .A(n113), .Y(n215) );
  CLKINVX1 U531 ( .A(n108), .Y(n214) );
  NAND2BX1 U532 ( .AN(n82), .B(n83), .Y(n10) );
  NAND2BX1 U533 ( .AN(n90), .B(n91), .Y(n12) );
  NAND2BX1 U534 ( .AN(n40), .B(n41), .Y(n3) );
  NAND2BX1 U535 ( .AN(n52), .B(n53), .Y(n5) );
  NAND2X1 U536 ( .A(n372), .B(n38), .Y(n2) );
  NAND2BX1 U537 ( .AN(n100), .B(n101), .Y(n13) );
  NAND2BX1 U538 ( .AN(n87), .B(n88), .Y(n11) );
  NAND2BX1 U539 ( .AN(n79), .B(n80), .Y(n9) );
  NAND2BX1 U540 ( .AN(n66), .B(n67), .Y(n7) );
  CLKINVX1 U541 ( .A(n185), .Y(n183) );
  CLKINVX1 U542 ( .A(n154), .Y(n152) );
  NAND2X1 U543 ( .A(n230), .B(n198), .Y(n31) );
  NAND2X1 U544 ( .A(n229), .B(n194), .Y(n30) );
  CLKINVX1 U545 ( .A(n193), .Y(n229) );
  INVXL U546 ( .A(B[12]), .Y(n250) );
  INVXL U547 ( .A(B[10]), .Y(n252) );
  INVXL U548 ( .A(B[11]), .Y(n251) );
  INVXL U549 ( .A(B[9]), .Y(n253) );
  INVXL U550 ( .A(B[6]), .Y(n256) );
  INVXL U551 ( .A(B[14]), .Y(n248) );
  INVXL U552 ( .A(B[15]), .Y(n247) );
  INVXL U553 ( .A(B[5]), .Y(n257) );
  INVXL U554 ( .A(B[3]), .Y(n259) );
  INVXL U555 ( .A(B[4]), .Y(n258) );
  NOR2X1 U556 ( .A(n259), .B(A[3]), .Y(n190) );
  NOR2X1 U557 ( .A(n256), .B(A[6]), .Y(n174) );
  NOR2X1 U558 ( .A(n257), .B(A[5]), .Y(n179) );
  NAND2X1 U559 ( .A(n248), .B(A[14]), .Y(n129) );
  NAND2X1 U560 ( .A(n256), .B(A[6]), .Y(n175) );
  NAND2X1 U561 ( .A(n244), .B(A[18]), .Y(n104) );
  NAND2X1 U562 ( .A(n250), .B(A[12]), .Y(n141) );
  NAND2X1 U563 ( .A(n246), .B(A[16]), .Y(n114) );
  NOR2X1 U564 ( .A(n248), .B(A[14]), .Y(n128) );
  NOR2X1 U565 ( .A(n250), .B(A[12]), .Y(n140) );
  NOR2X1 U566 ( .A(n252), .B(A[10]), .Y(n153) );
  NOR2X1 U567 ( .A(n261), .B(A[1]), .Y(n197) );
  NOR2X1 U568 ( .A(n262), .B(A[0]), .Y(n199) );
  NOR2X1 U569 ( .A(n238), .B(A[24]), .Y(n69) );
  OR2X1 U570 ( .A(n236), .B(A[26]), .Y(n371) );
  OR2X1 U571 ( .A(n32), .B(n374), .Y(n1) );
endmodule


module Execution_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n34, n37, n39, n40, n41, n42, n43, n45, n47, n48, n49, n50, n51,
         n52, n53, n54, n55, n56, n57, n58, n59, n61, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n201,
         n204, n206, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n337, n338, n339, n340, n341, n342,
         n343, n344, n345;

  AOI21XL U269 ( .A0(n87), .A1(n78), .B0(n79), .Y(n77) );
  OAI21X1 U270 ( .A0(n88), .A1(n92), .B0(n89), .Y(n87) );
  NAND2XL U271 ( .A(n229), .B(n186), .Y(n28) );
  INVXL U272 ( .A(n186), .Y(n184) );
  OAI21X2 U273 ( .A0(n180), .A1(n186), .B0(n181), .Y(n179) );
  NOR2X6 U274 ( .A(B[3]), .B(A[3]), .Y(n191) );
  NAND2X4 U275 ( .A(B[3]), .B(A[3]), .Y(n192) );
  NOR2X1 U276 ( .A(B[6]), .B(A[6]), .Y(n175) );
  NAND2X1 U277 ( .A(B[6]), .B(A[6]), .Y(n176) );
  NOR2X1 U278 ( .A(n80), .B(n83), .Y(n78) );
  AOI21X1 U279 ( .A0(n197), .A1(n189), .B0(n190), .Y(n188) );
  OAI21XL U280 ( .A0(n191), .A1(n195), .B0(n192), .Y(n190) );
  OAI21XL U281 ( .A0(n149), .A1(n155), .B0(n150), .Y(n148) );
  NOR2X1 U282 ( .A(B[17]), .B(A[17]), .Y(n109) );
  OAI21XL U283 ( .A0(n59), .A1(n53), .B0(n54), .Y(n52) );
  NOR2X1 U284 ( .A(B[1]), .B(A[1]), .Y(n198) );
  NOR2X1 U285 ( .A(B[7]), .B(A[7]), .Y(n172) );
  NOR2X1 U286 ( .A(B[19]), .B(A[19]), .Y(n101) );
  OAI21XL U287 ( .A0(n109), .A1(n115), .B0(n110), .Y(n108) );
  NOR2X1 U288 ( .A(B[23]), .B(A[23]), .Y(n80) );
  NOR2X1 U289 ( .A(n70), .B(n67), .Y(n65) );
  NOR2X1 U290 ( .A(n88), .B(n91), .Y(n86) );
  NOR2X1 U291 ( .A(B[27]), .B(A[27]), .Y(n53) );
  NOR2X1 U292 ( .A(n337), .B(n75), .Y(n73) );
  NAND2X1 U293 ( .A(B[2]), .B(A[2]), .Y(n195) );
  OAI21X1 U294 ( .A0(n143), .A1(n132), .B0(n133), .Y(n131) );
  NOR2X1 U295 ( .A(B[21]), .B(A[21]), .Y(n88) );
  NOR2X1 U296 ( .A(B[20]), .B(A[20]), .Y(n91) );
  NAND2X1 U297 ( .A(B[18]), .B(A[18]), .Y(n105) );
  OR2X1 U298 ( .A(B[26]), .B(A[26]), .Y(n341) );
  NOR2X1 U299 ( .A(B[22]), .B(A[22]), .Y(n83) );
  AND2X2 U300 ( .A(n344), .B(n201), .Y(SUM[0]) );
  NAND2X1 U301 ( .A(B[12]), .B(A[12]), .Y(n142) );
  INVX3 U302 ( .A(n117), .Y(n116) );
  NAND2X1 U303 ( .A(B[16]), .B(A[16]), .Y(n115) );
  NOR2X1 U304 ( .A(B[13]), .B(A[13]), .Y(n136) );
  NOR2X1 U305 ( .A(B[18]), .B(A[18]), .Y(n104) );
  NOR2XL U306 ( .A(B[16]), .B(A[16]), .Y(n114) );
  NAND2XL U307 ( .A(B[13]), .B(A[13]), .Y(n137) );
  NAND2X1 U308 ( .A(B[0]), .B(A[0]), .Y(n201) );
  NAND2XL U309 ( .A(B[1]), .B(A[1]), .Y(n199) );
  CLKINVX1 U310 ( .A(n73), .Y(n72) );
  OAI21XL U311 ( .A0(n80), .A1(n84), .B0(n81), .Y(n79) );
  OAI21XL U312 ( .A0(n73), .A1(n70), .B0(n71), .Y(n69) );
  NOR2X1 U313 ( .A(B[25]), .B(A[25]), .Y(n67) );
  AND2XL U314 ( .A(n116), .B(n74), .Y(n337) );
  OAI21X2 U315 ( .A0(n98), .A1(n76), .B0(n77), .Y(n75) );
  NOR2X1 U316 ( .A(n76), .B(n97), .Y(n74) );
  NAND2X2 U317 ( .A(n134), .B(n122), .Y(n120) );
  INVXL U318 ( .A(n87), .Y(n339) );
  NOR2XL U319 ( .A(n164), .B(n161), .Y(n159) );
  NAND2XL U320 ( .A(n220), .B(n137), .Y(n19) );
  INVXL U321 ( .A(n136), .Y(n220) );
  INVXL U322 ( .A(n91), .Y(n213) );
  NOR2X1 U323 ( .A(B[14]), .B(A[14]), .Y(n129) );
  NAND2XL U324 ( .A(B[4]), .B(A[4]), .Y(n186) );
  NAND2XL U325 ( .A(B[19]), .B(A[19]), .Y(n102) );
  NAND2X2 U326 ( .A(B[8]), .B(A[8]), .Y(n165) );
  NOR2X2 U327 ( .A(B[8]), .B(A[8]), .Y(n164) );
  INVX3 U328 ( .A(n94), .Y(n93) );
  OAI21X1 U329 ( .A0(n146), .A1(n120), .B0(n121), .Y(n119) );
  NAND2X1 U330 ( .A(n159), .B(n147), .Y(n145) );
  INVXL U331 ( .A(n59), .Y(n57) );
  INVXL U332 ( .A(n197), .Y(n196) );
  NAND2X1 U333 ( .A(n93), .B(n86), .Y(n338) );
  AND2X2 U334 ( .A(n338), .B(n339), .Y(n85) );
  AOI21X1 U335 ( .A0(n135), .A1(n122), .B0(n123), .Y(n121) );
  NOR2X1 U336 ( .A(n129), .B(n124), .Y(n122) );
  OAI21X1 U337 ( .A0(n136), .A1(n142), .B0(n137), .Y(n135) );
  OAI21XL U338 ( .A0(n106), .A1(n104), .B0(n105), .Y(n103) );
  OAI21X1 U339 ( .A0(n43), .A1(n41), .B0(n42), .Y(n40) );
  NOR2X1 U340 ( .A(n141), .B(n136), .Y(n134) );
  OAI21X1 U341 ( .A0(n67), .A1(n71), .B0(n68), .Y(n66) );
  INVXL U342 ( .A(n198), .Y(n232) );
  OAI21XL U343 ( .A0(n85), .A1(n83), .B0(n84), .Y(n82) );
  XOR2X1 U344 ( .A(n85), .B(n10), .Y(SUM[22]) );
  INVXL U345 ( .A(n58), .Y(n56) );
  OAI21XL U346 ( .A0(n166), .A1(n145), .B0(n146), .Y(n144) );
  AOI21XL U347 ( .A0(n187), .A1(n178), .B0(n179), .Y(n177) );
  AOI21XL U348 ( .A0(n116), .A1(n107), .B0(n108), .Y(n106) );
  INVX1 U349 ( .A(n167), .Y(n166) );
  NAND2XL U350 ( .A(n224), .B(n162), .Y(n23) );
  INVXL U351 ( .A(n161), .Y(n224) );
  NAND2XL U352 ( .A(n226), .B(n173), .Y(n25) );
  INVXL U353 ( .A(n172), .Y(n226) );
  NAND2XL U354 ( .A(n211), .B(n84), .Y(n10) );
  INVXL U355 ( .A(n83), .Y(n211) );
  XOR2XL U356 ( .A(n143), .B(n20), .Y(SUM[12]) );
  INVXL U357 ( .A(n88), .Y(n212) );
  AOI21XL U358 ( .A0(n116), .A1(n217), .B0(n113), .Y(n111) );
  NAND2XL U359 ( .A(n222), .B(n150), .Y(n21) );
  INVXL U360 ( .A(n149), .Y(n222) );
  AOI21XL U361 ( .A0(n144), .A1(n221), .B0(n140), .Y(n138) );
  NAND2XL U362 ( .A(n218), .B(n125), .Y(n17) );
  INVXL U363 ( .A(n124), .Y(n218) );
  NAND2XL U364 ( .A(n230), .B(n192), .Y(n29) );
  INVXL U365 ( .A(n191), .Y(n230) );
  NAND2XL U366 ( .A(n232), .B(n199), .Y(n31) );
  NAND2XL U367 ( .A(n228), .B(n181), .Y(n27) );
  AOI21XL U368 ( .A0(n187), .A1(n229), .B0(n184), .Y(n182) );
  INVXL U369 ( .A(n180), .Y(n228) );
  XOR2XL U370 ( .A(n166), .B(n24), .Y(SUM[8]) );
  INVXL U371 ( .A(n164), .Y(n225) );
  XOR2XL U372 ( .A(n196), .B(n30), .Y(SUM[2]) );
  INVXL U373 ( .A(n194), .Y(n231) );
  XOR2XL U374 ( .A(n177), .B(n26), .Y(SUM[6]) );
  INVXL U375 ( .A(n175), .Y(n227) );
  XNOR2XL U376 ( .A(n187), .B(n28), .Y(SUM[4]) );
  INVXL U377 ( .A(n70), .Y(n209) );
  INVXL U378 ( .A(n109), .Y(n216) );
  INVXL U379 ( .A(n80), .Y(n210) );
  INVXL U380 ( .A(n101), .Y(n214) );
  INVXL U381 ( .A(n53), .Y(n206) );
  NAND2XL U382 ( .A(B[10]), .B(A[10]), .Y(n155) );
  NOR2XL U383 ( .A(B[12]), .B(A[12]), .Y(n141) );
  NAND2XL U384 ( .A(B[14]), .B(A[14]), .Y(n130) );
  XNOR2X1 U385 ( .A(n340), .B(n1), .Y(SUM[31]) );
  AO21X1 U386 ( .A0(n40), .A1(n342), .B0(n37), .Y(n340) );
  NOR2XL U387 ( .A(B[10]), .B(A[10]), .Y(n154) );
  NOR2XL U388 ( .A(B[4]), .B(A[4]), .Y(n185) );
  NAND2XL U389 ( .A(B[21]), .B(A[21]), .Y(n89) );
  NAND2XL U390 ( .A(B[26]), .B(A[26]), .Y(n63) );
  NAND2XL U391 ( .A(B[23]), .B(A[23]), .Y(n81) );
  NAND2XL U392 ( .A(B[27]), .B(A[27]), .Y(n54) );
  NOR2XL U393 ( .A(B[29]), .B(A[29]), .Y(n41) );
  NAND2XL U394 ( .A(B[30]), .B(A[30]), .Y(n39) );
  NAND2XL U395 ( .A(B[29]), .B(A[29]), .Y(n42) );
  OR2XL U396 ( .A(B[30]), .B(A[30]), .Y(n342) );
  OR2XL U397 ( .A(B[31]), .B(A[31]), .Y(n345) );
  OR2XL U398 ( .A(B[0]), .B(A[0]), .Y(n344) );
  CLKINVX1 U399 ( .A(n144), .Y(n143) );
  AOI21X1 U400 ( .A0(n116), .A1(n95), .B0(n96), .Y(n94) );
  CLKINVX1 U401 ( .A(n97), .Y(n95) );
  CLKINVX1 U402 ( .A(n98), .Y(n96) );
  AOI21X1 U403 ( .A0(n167), .A1(n118), .B0(n119), .Y(n117) );
  NOR2X1 U404 ( .A(n145), .B(n120), .Y(n118) );
  OAI21XL U405 ( .A0(n166), .A1(n157), .B0(n158), .Y(n156) );
  CLKINVX1 U406 ( .A(n159), .Y(n157) );
  CLKINVX1 U407 ( .A(n160), .Y(n158) );
  CLKINVX1 U408 ( .A(n134), .Y(n132) );
  CLKINVX1 U409 ( .A(n135), .Y(n133) );
  AOI21X1 U410 ( .A0(n72), .A1(n65), .B0(n66), .Y(n64) );
  AOI21X1 U411 ( .A0(n72), .A1(n56), .B0(n57), .Y(n55) );
  CLKINVX1 U412 ( .A(n188), .Y(n187) );
  NAND2X1 U413 ( .A(n78), .B(n86), .Y(n76) );
  XOR2X1 U414 ( .A(n64), .B(n6), .Y(SUM[26]) );
  NAND2X1 U415 ( .A(n99), .B(n107), .Y(n97) );
  OAI21X1 U416 ( .A0(n161), .A1(n165), .B0(n162), .Y(n160) );
  OAI21X1 U417 ( .A0(n198), .A1(n201), .B0(n199), .Y(n197) );
  AOI21X1 U418 ( .A0(n48), .A1(n343), .B0(n45), .Y(n43) );
  CLKINVX1 U419 ( .A(n47), .Y(n45) );
  OAI21X1 U420 ( .A0(n188), .A1(n168), .B0(n169), .Y(n167) );
  NAND2X1 U421 ( .A(n170), .B(n178), .Y(n168) );
  AOI21X1 U422 ( .A0(n179), .A1(n170), .B0(n171), .Y(n169) );
  NOR2X1 U423 ( .A(n175), .B(n172), .Y(n170) );
  AOI21X1 U424 ( .A0(n66), .A1(n341), .B0(n61), .Y(n59) );
  CLKINVX1 U425 ( .A(n63), .Y(n61) );
  AOI21X1 U426 ( .A0(n108), .A1(n99), .B0(n100), .Y(n98) );
  OAI21XL U427 ( .A0(n101), .A1(n105), .B0(n102), .Y(n100) );
  NOR2X1 U428 ( .A(n194), .B(n191), .Y(n189) );
  AOI21X1 U429 ( .A0(n160), .A1(n147), .B0(n148), .Y(n146) );
  OAI21X1 U430 ( .A0(n117), .A1(n49), .B0(n50), .Y(n48) );
  NAND2X1 U431 ( .A(n51), .B(n74), .Y(n49) );
  AOI21X1 U432 ( .A0(n75), .A1(n51), .B0(n52), .Y(n50) );
  NOR2X1 U433 ( .A(n58), .B(n53), .Y(n51) );
  XNOR2X1 U434 ( .A(n90), .B(n11), .Y(SUM[21]) );
  NAND2X1 U435 ( .A(n212), .B(n89), .Y(n11) );
  OAI21XL U436 ( .A0(n94), .A1(n91), .B0(n92), .Y(n90) );
  XNOR2X1 U437 ( .A(n156), .B(n22), .Y(SUM[10]) );
  NAND2X1 U438 ( .A(n223), .B(n155), .Y(n22) );
  XNOR2X1 U439 ( .A(n131), .B(n18), .Y(SUM[14]) );
  NAND2X1 U440 ( .A(n219), .B(n130), .Y(n18) );
  XNOR2X1 U441 ( .A(n163), .B(n23), .Y(SUM[9]) );
  OAI21XL U442 ( .A0(n166), .A1(n164), .B0(n165), .Y(n163) );
  XNOR2X1 U443 ( .A(n174), .B(n25), .Y(SUM[7]) );
  OAI21XL U444 ( .A0(n177), .A1(n175), .B0(n176), .Y(n174) );
  OAI21XL U445 ( .A0(n172), .A1(n176), .B0(n173), .Y(n171) );
  NOR2X1 U446 ( .A(n180), .B(n185), .Y(n178) );
  NOR2X1 U447 ( .A(n154), .B(n149), .Y(n147) );
  NOR2X1 U448 ( .A(n101), .B(n104), .Y(n99) );
  CLKINVX1 U449 ( .A(n115), .Y(n113) );
  OAI21XL U450 ( .A0(n124), .A1(n130), .B0(n125), .Y(n123) );
  XOR2X1 U451 ( .A(n55), .B(n5), .Y(SUM[27]) );
  NAND2X1 U452 ( .A(n206), .B(n54), .Y(n5) );
  XNOR2X1 U453 ( .A(n40), .B(n2), .Y(SUM[30]) );
  NAND2X1 U454 ( .A(n342), .B(n39), .Y(n2) );
  XOR2X1 U455 ( .A(n106), .B(n14), .Y(SUM[18]) );
  NAND2X1 U456 ( .A(n215), .B(n105), .Y(n14) );
  XNOR2X1 U457 ( .A(n116), .B(n16), .Y(SUM[16]) );
  NAND2X1 U458 ( .A(n217), .B(n115), .Y(n16) );
  XNOR2X1 U459 ( .A(n82), .B(n9), .Y(SUM[23]) );
  NAND2X1 U460 ( .A(n210), .B(n81), .Y(n9) );
  XNOR2X1 U461 ( .A(n93), .B(n12), .Y(SUM[20]) );
  NAND2X1 U462 ( .A(n213), .B(n92), .Y(n12) );
  XOR2X1 U463 ( .A(n111), .B(n15), .Y(SUM[17]) );
  NAND2X1 U464 ( .A(n216), .B(n110), .Y(n15) );
  XNOR2X1 U465 ( .A(n103), .B(n13), .Y(SUM[19]) );
  NAND2X1 U466 ( .A(n214), .B(n102), .Y(n13) );
  XNOR2X1 U467 ( .A(n48), .B(n4), .Y(SUM[28]) );
  NAND2X1 U468 ( .A(n343), .B(n47), .Y(n4) );
  XNOR2X1 U469 ( .A(n72), .B(n8), .Y(SUM[24]) );
  NAND2X1 U470 ( .A(n209), .B(n71), .Y(n8) );
  XOR2X1 U471 ( .A(n43), .B(n3), .Y(SUM[29]) );
  NAND2X1 U472 ( .A(n204), .B(n42), .Y(n3) );
  XNOR2X1 U473 ( .A(n69), .B(n7), .Y(SUM[25]) );
  NAND2X1 U474 ( .A(n208), .B(n68), .Y(n7) );
  XOR2X1 U475 ( .A(n182), .B(n27), .Y(SUM[5]) );
  XOR2X1 U476 ( .A(n126), .B(n17), .Y(SUM[15]) );
  AOI21X1 U477 ( .A0(n131), .A1(n219), .B0(n128), .Y(n126) );
  NAND2X1 U478 ( .A(n221), .B(n142), .Y(n20) );
  XOR2X1 U479 ( .A(n151), .B(n21), .Y(SUM[11]) );
  AOI21X1 U480 ( .A0(n156), .A1(n223), .B0(n153), .Y(n151) );
  XOR2X1 U481 ( .A(n138), .B(n19), .Y(SUM[13]) );
  NAND2X1 U482 ( .A(n227), .B(n176), .Y(n26) );
  NAND2X1 U483 ( .A(n225), .B(n165), .Y(n24) );
  XNOR2X1 U484 ( .A(n193), .B(n29), .Y(SUM[3]) );
  OAI21XL U485 ( .A0(n196), .A1(n194), .B0(n195), .Y(n193) );
  NOR2X1 U486 ( .A(n109), .B(n114), .Y(n107) );
  CLKINVX1 U487 ( .A(n141), .Y(n221) );
  CLKINVX1 U488 ( .A(n154), .Y(n223) );
  CLKINVX1 U489 ( .A(n129), .Y(n219) );
  CLKINVX1 U490 ( .A(n185), .Y(n229) );
  CLKINVX1 U491 ( .A(n114), .Y(n217) );
  NAND2X1 U492 ( .A(n65), .B(n341), .Y(n58) );
  CLKINVX1 U493 ( .A(n104), .Y(n215) );
  CLKINVX1 U494 ( .A(n67), .Y(n208) );
  CLKINVX1 U495 ( .A(n142), .Y(n140) );
  CLKINVX1 U496 ( .A(n155), .Y(n153) );
  CLKINVX1 U497 ( .A(n130), .Y(n128) );
  CLKINVX1 U498 ( .A(n41), .Y(n204) );
  NAND2X1 U499 ( .A(n341), .B(n63), .Y(n6) );
  CLKINVX1 U500 ( .A(n39), .Y(n37) );
  XOR2X1 U501 ( .A(n31), .B(n201), .Y(SUM[1]) );
  NAND2X1 U502 ( .A(n231), .B(n195), .Y(n30) );
  NOR2X1 U503 ( .A(B[11]), .B(A[11]), .Y(n149) );
  NOR2X1 U504 ( .A(B[9]), .B(A[9]), .Y(n161) );
  NOR2X1 U505 ( .A(B[15]), .B(A[15]), .Y(n124) );
  NOR2X1 U506 ( .A(B[5]), .B(A[5]), .Y(n180) );
  NOR2X1 U507 ( .A(B[2]), .B(A[2]), .Y(n194) );
  NAND2XL U508 ( .A(B[11]), .B(A[11]), .Y(n150) );
  NAND2XL U509 ( .A(B[9]), .B(A[9]), .Y(n162) );
  NAND2XL U510 ( .A(B[15]), .B(A[15]), .Y(n125) );
  NAND2XL U511 ( .A(B[7]), .B(A[7]), .Y(n173) );
  NAND2XL U512 ( .A(B[5]), .B(A[5]), .Y(n181) );
  NAND2X1 U513 ( .A(B[24]), .B(A[24]), .Y(n71) );
  NAND2X1 U514 ( .A(B[20]), .B(A[20]), .Y(n92) );
  NAND2X1 U515 ( .A(B[17]), .B(A[17]), .Y(n110) );
  NAND2X1 U516 ( .A(B[25]), .B(A[25]), .Y(n68) );
  NAND2X1 U517 ( .A(n345), .B(n34), .Y(n1) );
  NAND2X1 U518 ( .A(B[31]), .B(A[31]), .Y(n34) );
  NOR2X1 U519 ( .A(B[24]), .B(A[24]), .Y(n70) );
  NAND2X1 U520 ( .A(B[22]), .B(A[22]), .Y(n84) );
  NAND2X1 U521 ( .A(B[28]), .B(A[28]), .Y(n47) );
  OR2X1 U522 ( .A(B[28]), .B(A[28]), .Y(n343) );
endmodule


module Execution_test_1 ( clk, rst, stall, ID_WB, ID_MEM, ID_EX, RData1, 
        RData2, Immediate_SE, ID_RegisterRt, ID_RegisterRd, WB, MEM, 
        next_ALUresult, ALUresult, MEMWriteData, RegisterRd, WBData, ForwardA, 
        ForwardB, test_si, test_so, test_se );
  input [1:0] ID_WB;
  input [2:0] ID_MEM;
  input [6:0] ID_EX;
  input [31:0] RData1;
  input [31:0] RData2;
  input [31:0] Immediate_SE;
  input [4:0] ID_RegisterRt;
  input [4:0] ID_RegisterRd;
  output [1:0] WB;
  output [2:0] MEM;
  output [31:0] next_ALUresult;
  output [31:0] ALUresult;
  output [31:0] MEMWriteData;
  output [4:0] RegisterRd;
  input [31:0] WBData;
  input [1:0] ForwardA;
  input [1:0] ForwardB;
  input clk, rst, stall, test_si, test_se;
  output test_so;
  wire   n1189, n1190, n1191, n1192, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, N172, N173, N174, N175, N176, N177, N178, N179, N180,
         N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191,
         N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202,
         N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213,
         N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224,
         N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235,
         N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342,
         N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353,
         N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N364,
         N365, N366, N367, N368, N369, N370, N371, N372, N373, N374, N375,
         N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386,
         N387, N388, N389, N390, N391, N392, N393, N394, N395, N493, N494,
         N495, N496, N497, N498, N499, N500, N501, N502, N503, N504, N505,
         N506, N507, N508, N524, n106, n129, n130, n139, n140, n156, n157,
         n158, n168, n177, n185, n186, n197, n198, n214, n215, n220, n231,
         n232, n247, n248, n268, n269, n295, n312, n313, n329, n330, n331,
         n348, n349, n350, n351, n353, n354, n358, n359, n428, n429, n431,
         n433, n434, n435, n439, n441, n442, n443, n444, n445, n446, n447,
         n448, n451, n453, n454, n455, n458, n461, n464, n467, n470, n473,
         n476, n479, n482, n485, n488, n491, n494, n497, n500, n503, n506,
         n509, n512, n515, n518, n521, n527, n530, n533, n536, n539, n542,
         n545, n549, n632, n633, n634, n635, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n61, n63, n65, n67, n69, n71, n73, n75, n77, n79, n1131, n99,
         n100, n101, n102, n103, n105, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n131, n132, n133, n134, n135, n136,
         n137, n138, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n169, n170, n171, n172, n173, n174, n175,
         n176, n178, n179, n180, n181, n182, n183, n184, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n216, n217, n218, n219, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n352, n355,
         n356, n357, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n430, n432, n436, n437, n438, n440, n449,
         n450, n452, n456, n457, n459, n460, n462, n463, n465, n466, n468,
         n469, n471, n472, n474, n475, n477, n478, n480, n481, n483, n484,
         n486, n487, n489, n490, n492, n493, n495, n496, n498, n499, n501,
         n502, n504, n505, n507, n508, n510, n511, n513, n514, n516, n517,
         n519, n520, n522, n523, n524, n525, n526, n528, n529, n531, n532,
         n534, n535, n537, n538, n540, n541, n543, n544, n546, n547, n548,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n636, n674, n675, n676, n677, n678,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1129, n3, n4, n36, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n62, n64, n66, n68, n70, n72, n74, n76, n78, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n104, n751, n764, n777, n791, n804, n817, n842, n855, n868, n892,
         n905, n950, n1041, n1130, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1146, n1147, n1148,
         n1149, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187;
  wire   [31:0] ALUData1;
  wire   [31:0] ALUData2;

  BUFX2 U3 ( .A(ALUData2[14]), .Y(n108) );
  BUFX4 U4 ( .A(n275), .Y(n277) );
  BUFX8 U5 ( .A(ALUData2[0]), .Y(n5) );
  OAI221XL U6 ( .A0(n1148), .A1(n283), .B0(n250), .B1(n1120), .C0(n934), .Y(
        ALUData2[0]) );
  BUFX6 U11 ( .A(n135), .Y(n6) );
  AND2XL U12 ( .A(n362), .B(n361), .Y(n135) );
  OAI221X2 U13 ( .A0(n1060), .A1(n281), .B0(n1095), .B1(n280), .C0(n750), .Y(
        ALUData2[14]) );
  BUFX16 U14 ( .A(n278), .Y(n280) );
  OAI221X4 U15 ( .A0(n1154), .A1(n276), .B0(n1071), .B1(n274), .C0(n890), .Y(
        ALUData1[3]) );
  NAND2X2 U16 ( .A(n352), .B(n357), .Y(n932) );
  OR2X4 U17 ( .A(ID_EX[0]), .B(ForwardB[1]), .Y(n356) );
  CLKBUFX3 U18 ( .A(ALUData2[30]), .Y(n252) );
  CLKBUFX3 U19 ( .A(ALUData2[28]), .Y(n254) );
  CLKBUFX3 U20 ( .A(ALUData2[21]), .Y(n264) );
  CLKBUFX3 U21 ( .A(ALUData2[19]), .Y(n266) );
  CLKBUFX3 U22 ( .A(ALUData2[18]), .Y(n267) );
  CLKBUFX3 U23 ( .A(ALUData2[23]), .Y(n262) );
  INVX1 U24 ( .A(n260), .Y(n725) );
  CLKBUFX3 U25 ( .A(ALUData2[22]), .Y(n263) );
  CLKBUFX3 U26 ( .A(ALUData2[27]), .Y(n255) );
  CLKINVX1 U27 ( .A(n995), .Y(n980) );
  CLKBUFX3 U28 ( .A(ALUData2[26]), .Y(n259) );
  CLKBUFX3 U29 ( .A(n998), .Y(n257) );
  NAND2XL U30 ( .A(RData1[24]), .B(n6), .Y(n426) );
  INVX1 U31 ( .A(n261), .Y(n724) );
  OR3X4 U32 ( .A(n99), .B(n100), .C(n101), .Y(ALUData2[13]) );
  CLKINVX1 U33 ( .A(n763), .Y(n101) );
  CLKINVX1 U34 ( .A(ForwardA[0]), .Y(n361) );
  CLKINVX1 U35 ( .A(ForwardA[1]), .Y(n362) );
  OAI221X1 U36 ( .A0(n1063), .A1(n281), .B0(n1098), .B1(n280), .C0(n790), .Y(
        ALUData2[11]) );
  CLKINVX1 U37 ( .A(Immediate_SE[9]), .Y(n316) );
  OR2X1 U38 ( .A(n312), .B(n313), .Y(n295) );
  NOR3X1 U39 ( .A(n317), .B(n315), .C(n308), .Y(n358) );
  NOR3X1 U40 ( .A(n307), .B(n315), .C(n317), .Y(n359) );
  CLKINVX1 U41 ( .A(Immediate_SE[10]), .Y(n318) );
  CLKBUFX6 U42 ( .A(n936), .Y(n283) );
  CLKINVX1 U43 ( .A(Immediate_SE[6]), .Y(n308) );
  CLKINVX1 U44 ( .A(Immediate_SE[7]), .Y(n310) );
  OR3X4 U45 ( .A(n105), .B(n107), .C(n7), .Y(ALUData2[8]) );
  MXI3X1 U46 ( .A(n235), .B(n236), .C(n193), .S0(n249), .S1(n246), .Y(n192) );
  CLKINVX1 U47 ( .A(n262), .Y(n621) );
  CLKBUFX3 U48 ( .A(ALUData2[29]), .Y(n253) );
  CLKINVX1 U49 ( .A(n255), .Y(n728) );
  CLKINVX1 U50 ( .A(WBData[3]), .Y(n1071) );
  CLKINVX1 U51 ( .A(WBData[8]), .Y(n1066) );
  CLKINVX1 U52 ( .A(WBData[12]), .Y(n1062) );
  CLKINVX1 U53 ( .A(WBData[15]), .Y(n1059) );
  AO22X1 U54 ( .A0(N179), .A1(n148), .B0(N371), .B1(n150), .Y(n849) );
  NAND4BX1 U55 ( .AN(n1007), .B(n1006), .C(n1005), .D(n1004), .Y(
        next_ALUresult[30]) );
  NAND4BX1 U56 ( .AN(n718), .B(n717), .C(n716), .D(n715), .Y(
        next_ALUresult[17]) );
  NAND4BX1 U57 ( .AN(n569), .B(n568), .C(n567), .D(n566), .Y(
        next_ALUresult[20]) );
  NAND4BX1 U58 ( .AN(n551), .B(n550), .C(n548), .D(n547), .Y(
        next_ALUresult[21]) );
  AOI221XL U59 ( .A0(N385), .A1(n150), .B0(N193), .B1(n148), .C0(n546), .Y(
        n547) );
  NAND4X1 U60 ( .A(n113), .B(n949), .C(n948), .D(n947), .Y(next_ALUresult[0])
         );
  NAND4X1 U61 ( .A(n110), .B(n960), .C(n959), .D(n958), .Y(next_ALUresult[15])
         );
  NAND4X1 U62 ( .A(n115), .B(n787), .C(n786), .D(n785), .Y(next_ALUresult[12])
         );
  NAND4BX1 U63 ( .AN(n590), .B(n589), .C(n588), .D(n587), .Y(
        next_ALUresult[19]) );
  NAND4BX1 U64 ( .AN(n614), .B(n613), .C(n612), .D(n611), .Y(
        next_ALUresult[18]) );
  NAND4BX2 U65 ( .AN(n492), .B(n490), .C(n489), .D(n487), .Y(
        next_ALUresult[23]) );
  NAND4BX1 U66 ( .AN(n408), .B(n407), .C(n406), .D(n405), .Y(
        next_ALUresult[26]) );
  CLKMX2X2 U67 ( .A(n1026), .B(ALUresult[31]), .S0(n320), .Y(
        next_ALUresult[31]) );
  NAND3BX1 U68 ( .AN(n1025), .B(n1024), .C(n1023), .Y(n1026) );
  NAND4BX1 U69 ( .AN(n425), .B(n424), .C(n423), .D(n422), .Y(
        next_ALUresult[25]) );
  NAND4BX2 U70 ( .AN(n520), .B(n519), .C(n517), .D(n516), .Y(
        next_ALUresult[22]) );
  AOI221XL U71 ( .A0(N386), .A1(n150), .B0(N194), .B1(n298), .C0(n514), .Y(
        n516) );
  NAND4BX1 U72 ( .AN(n393), .B(n392), .C(n391), .D(n390), .Y(
        next_ALUresult[27]) );
  NAND4BX1 U73 ( .AN(n465), .B(n463), .C(n462), .D(n460), .Y(
        next_ALUresult[24]) );
  NAND4X1 U74 ( .A(n119), .B(n774), .C(n773), .D(n772), .Y(next_ALUresult[13])
         );
  NAND4X1 U75 ( .A(n112), .B(n801), .C(n800), .D(n799), .Y(next_ALUresult[11])
         );
  NAND4X1 U76 ( .A(n111), .B(n761), .C(n760), .D(n759), .Y(next_ALUresult[14])
         );
  CLKBUFX2 U77 ( .A(n932), .Y(n279) );
  CLKINVX1 U78 ( .A(ALUData2[4]), .Y(n235) );
  CLKBUFX6 U79 ( .A(n272), .Y(n273) );
  CLKINVX1 U80 ( .A(ALUData2[3]), .Y(n896) );
  CLKINVX1 U81 ( .A(ALUData2[2]), .Y(n234) );
  NAND2X1 U82 ( .A(n357), .B(n356), .Y(n936) );
  INVX4 U83 ( .A(n250), .Y(n789) );
  OAI22XL U84 ( .A0(n1066), .A1(n282), .B0(n1101), .B1(n280), .Y(n7) );
  CLKBUFX3 U85 ( .A(ALUData2[31]), .Y(n251) );
  NAND3X2 U86 ( .A(n102), .B(n103), .C(n916), .Y(ALUData2[1]) );
  CLKINVX1 U87 ( .A(ID_EX[0]), .Y(n347) );
  MXI2X1 U88 ( .A(n208), .B(n207), .S0(n246), .Y(n8) );
  MXI2X1 U89 ( .A(n212), .B(n211), .S0(n246), .Y(n9) );
  MXI2X1 U90 ( .A(n218), .B(n217), .S0(n246), .Y(n10) );
  CLKINVX1 U91 ( .A(ALUData2[5]), .Y(n236) );
  CLKINVX1 U92 ( .A(Immediate_SE[2]), .Y(n1118) );
  CLKINVX1 U93 ( .A(Immediate_SE[1]), .Y(n1119) );
  CLKINVX1 U94 ( .A(Immediate_SE[0]), .Y(n1120) );
  CLKINVX1 U95 ( .A(n535), .Y(n997) );
  NAND2X1 U96 ( .A(n348), .B(n359), .Y(n186) );
  INVX3 U97 ( .A(n308), .Y(n307) );
  INVX12 U98 ( .A(n26), .Y(MEMWriteData[16]) );
  INVX12 U99 ( .A(n25), .Y(MEMWriteData[20]) );
  INVX12 U100 ( .A(n24), .Y(MEMWriteData[18]) );
  INVX12 U101 ( .A(n23), .Y(MEMWriteData[17]) );
  INVX12 U102 ( .A(n35), .Y(MEMWriteData[2]) );
  INVX12 U103 ( .A(n34), .Y(MEMWriteData[3]) );
  INVX12 U104 ( .A(n33), .Y(MEMWriteData[4]) );
  INVX12 U105 ( .A(n32), .Y(MEMWriteData[5]) );
  INVX12 U106 ( .A(n31), .Y(MEMWriteData[6]) );
  INVX12 U107 ( .A(n30), .Y(MEMWriteData[7]) );
  INVX12 U108 ( .A(n29), .Y(MEMWriteData[8]) );
  INVX12 U109 ( .A(n28), .Y(MEMWriteData[9]) );
  INVX12 U110 ( .A(n27), .Y(MEMWriteData[10]) );
  INVX12 U111 ( .A(n22), .Y(MEMWriteData[11]) );
  INVX12 U112 ( .A(n21), .Y(MEMWriteData[12]) );
  INVX12 U113 ( .A(n20), .Y(MEMWriteData[13]) );
  INVX12 U114 ( .A(n19), .Y(MEMWriteData[14]) );
  INVX12 U115 ( .A(n18), .Y(MEMWriteData[15]) );
  INVX12 U116 ( .A(n17), .Y(MEMWriteData[26]) );
  INVX12 U117 ( .A(n16), .Y(MEMWriteData[25]) );
  INVX12 U118 ( .A(n15), .Y(MEMWriteData[24]) );
  INVX12 U119 ( .A(n14), .Y(MEMWriteData[23]) );
  INVX12 U120 ( .A(n13), .Y(MEMWriteData[22]) );
  INVX12 U121 ( .A(n12), .Y(MEMWriteData[21]) );
  INVX12 U122 ( .A(n11), .Y(MEMWriteData[19]) );
  CLKINVX1 U123 ( .A(n990), .Y(n61) );
  INVX16 U124 ( .A(n61), .Y(ALUresult[30]) );
  CLKINVX1 U125 ( .A(n617), .Y(n63) );
  INVX16 U126 ( .A(n63), .Y(ALUresult[17]) );
  CLKINVX1 U127 ( .A(n880), .Y(n65) );
  INVX16 U128 ( .A(n65), .Y(ALUresult[4]) );
  CLKINVX1 U129 ( .A(n721), .Y(n67) );
  INVX16 U130 ( .A(n67), .Y(ALUresult[16]) );
  CLKINVX1 U131 ( .A(n974), .Y(n69) );
  INVX16 U132 ( .A(n69), .Y(ALUresult[29]) );
  CLKINVX1 U133 ( .A(n961), .Y(n71) );
  INVX16 U134 ( .A(n71), .Y(ALUresult[28]) );
  CLKINVX1 U135 ( .A(n554), .Y(n73) );
  INVX16 U136 ( .A(n73), .Y(ALUresult[20]) );
  CLKINVX1 U137 ( .A(n524), .Y(n75) );
  INVX16 U138 ( .A(n75), .Y(ALUresult[21]) );
  CLKINVX1 U139 ( .A(n829), .Y(n77) );
  INVX16 U140 ( .A(n77), .Y(ALUresult[8]) );
  CLKINVX1 U141 ( .A(n917), .Y(n79) );
  INVX16 U142 ( .A(n79), .Y(ALUresult[1]) );
  OAI221X4 U143 ( .A0(n1175), .A1(n283), .B0(n250), .B1(n310), .C0(n841), .Y(
        ALUData2[7]) );
  OAI221X4 U144 ( .A0(n1187), .A1(n283), .B0(n250), .B1(n308), .C0(n854), .Y(
        ALUData2[6]) );
  OAI221X4 U145 ( .A0(n1178), .A1(n283), .B0(n250), .B1(n867), .C0(n866), .Y(
        ALUData2[5]) );
  OA22XL U146 ( .A0(n1069), .A1(n281), .B0(n1104), .B1(n279), .Y(n866) );
  OAI221X4 U147 ( .A0(n1153), .A1(n283), .B0(n250), .B1(n1117), .C0(n891), .Y(
        ALUData2[3]) );
  OA22XL U148 ( .A0(n1071), .A1(n282), .B0(n1106), .B1(n279), .Y(n891) );
  OAI221X4 U149 ( .A0(n1183), .A1(n283), .B0(n250), .B1(n1118), .C0(n904), .Y(
        ALUData2[2]) );
  OAI221X4 U150 ( .A0(n1059), .A1(n281), .B0(n1094), .B1(n280), .C0(n748), .Y(
        ALUData2[15]) );
  OAI221X4 U151 ( .A0(n1171), .A1(n283), .B0(n250), .B1(n316), .C0(n816), .Y(
        ALUData2[9]) );
  OA22XL U152 ( .A0(n1065), .A1(n282), .B0(n1100), .B1(n279), .Y(n816) );
  OAI221X4 U153 ( .A0(n1062), .A1(n281), .B0(n1097), .B1(n280), .C0(n776), .Y(
        ALUData2[12]) );
  OAI221X4 U154 ( .A0(n1181), .A1(n283), .B0(n250), .B1(n318), .C0(n803), .Y(
        ALUData2[10]) );
  OA22XL U155 ( .A0(n1064), .A1(n282), .B0(n1099), .B1(n278), .Y(n803) );
  INVX12 U156 ( .A(n892), .Y(MEMWriteData[0]) );
  INVX12 U157 ( .A(n1041), .Y(MEMWriteData[31]) );
  INVX12 U158 ( .A(n1133), .Y(MEMWriteData[30]) );
  INVX12 U159 ( .A(n1136), .Y(MEMWriteData[29]) );
  INVX12 U161 ( .A(n1139), .Y(MEMWriteData[28]) );
  INVX12 U162 ( .A(n1142), .Y(MEMWriteData[27]) );
  BUFX16 U163 ( .A(n1128), .Y(ALUresult[0]) );
  INVX16 U164 ( .A(n104), .Y(ALUresult[9]) );
  INVX16 U165 ( .A(n94), .Y(ALUresult[15]) );
  NAND4X1 U166 ( .A(n116), .B(n852), .C(n851), .D(n850), .Y(next_ALUresult[7])
         );
  INVX16 U167 ( .A(n751), .Y(ALUresult[7]) );
  INVX16 U168 ( .A(n95), .Y(ALUresult[12]) );
  BUFX16 U169 ( .A(n1126), .Y(ALUresult[19]) );
  BUFX16 U170 ( .A(n1127), .Y(ALUresult[18]) );
  NAND4X1 U171 ( .A(n123), .B(n889), .C(n888), .D(n887), .Y(next_ALUresult[4])
         );
  BUFX16 U172 ( .A(n1124), .Y(ALUresult[23]) );
  NAND4BX1 U173 ( .AN(n746), .B(n745), .C(n744), .D(n743), .Y(
        next_ALUresult[16]) );
  BUFX16 U174 ( .A(n1123), .Y(ALUresult[26]) );
  BUFX16 U175 ( .A(n1121), .Y(ALUresult[31]) );
  NAND4BX1 U176 ( .AN(n989), .B(n988), .C(n987), .D(n986), .Y(
        next_ALUresult[29]) );
  NAND4BX1 U177 ( .AN(n973), .B(n972), .C(n971), .D(n970), .Y(
        next_ALUresult[28]) );
  BUFX16 U178 ( .A(n411), .Y(ALUresult[25]) );
  INVX16 U179 ( .A(n764), .Y(ALUresult[5]) );
  BUFX16 U180 ( .A(n1125), .Y(ALUresult[22]) );
  BUFX16 U181 ( .A(n1122), .Y(ALUresult[27]) );
  BUFX16 U182 ( .A(n430), .Y(ALUresult[24]) );
  NAND4X1 U183 ( .A(n114), .B(n814), .C(n813), .D(n812), .Y(next_ALUresult[10]) );
  INVX16 U184 ( .A(n777), .Y(ALUresult[10]) );
  NAND4X1 U185 ( .A(n122), .B(n914), .C(n913), .D(n912), .Y(next_ALUresult[2])
         );
  INVX16 U186 ( .A(n791), .Y(ALUresult[2]) );
  NAND4X1 U187 ( .A(n121), .B(n902), .C(n901), .D(n900), .Y(next_ALUresult[3])
         );
  INVX16 U188 ( .A(n93), .Y(ALUresult[3]) );
  NAND4X1 U189 ( .A(n117), .B(n839), .C(n838), .D(n837), .Y(next_ALUresult[8])
         );
  NAND4X1 U190 ( .A(n118), .B(n864), .C(n863), .D(n862), .Y(next_ALUresult[6])
         );
  INVX16 U191 ( .A(n804), .Y(ALUresult[6]) );
  INVX16 U192 ( .A(n96), .Y(ALUresult[13]) );
  INVX16 U193 ( .A(n97), .Y(ALUresult[11]) );
  INVX16 U194 ( .A(n98), .Y(ALUresult[14]) );
  CLKINVX1 U195 ( .A(WBData[5]), .Y(n1069) );
  CLKINVX1 U196 ( .A(WBData[10]), .Y(n1064) );
  CLKINVX1 U197 ( .A(WBData[2]), .Y(n1072) );
  CLKINVX1 U198 ( .A(WBData[7]), .Y(n1067) );
  CLKINVX1 U199 ( .A(WBData[6]), .Y(n1068) );
  NAND2XL U200 ( .A(RData1[10]), .B(n6), .Y(n802) );
  MXI2X1 U201 ( .A(n144), .B(n137), .S0(Immediate_SE[8]), .Y(n184) );
  CLKBUFX3 U202 ( .A(n933), .Y(n281) );
  AOI2BB2XL U203 ( .B0(Immediate_SE[12]), .B1(n789), .A0N(n1159), .A1N(n283), 
        .Y(n776) );
  NAND2XL U204 ( .A(RData1[0]), .B(n6), .Y(n929) );
  OA22XL U205 ( .A0(n282), .A1(n1039), .B0(n278), .B1(n1040), .Y(n916) );
  OR2XL U206 ( .A(n710), .B(n283), .Y(n102) );
  OR2XL U207 ( .A(n250), .B(n1119), .Y(n103) );
  NOR2XL U208 ( .A(n1061), .B(n281), .Y(n99) );
  NOR2XL U209 ( .A(n1096), .B(n280), .Y(n100) );
  OAI222XL U210 ( .A0(n158), .A1(n724), .B0(n157), .B1(n725), .C0(n130), .C1(
        n621), .Y(n531) );
  AOI22X1 U211 ( .A0(N336), .A1(n287), .B0(N208), .B1(n152), .Y(n123) );
  AOI2BB2XL U212 ( .B0(Immediate_SE[13]), .B1(n789), .A0N(n1162), .A1N(n283), 
        .Y(n763) );
  MXI4X1 U213 ( .A(n226), .B(n224), .C(n225), .D(n1018), .S0(n245), .S1(n246), 
        .Y(n145) );
  AND2X2 U214 ( .A(n106), .B(n980), .Y(n109) );
  AO22X2 U215 ( .A0(N185), .A1(n298), .B0(N377), .B1(n297), .Y(n771) );
  MXI4X1 U216 ( .A(n204), .B(n209), .C(n210), .D(n1018), .S0(n245), .S1(n246), 
        .Y(n147) );
  MXI2X1 U217 ( .A(n191), .B(n187), .S0(Immediate_SE[7]), .Y(N498) );
  MXI4X1 U218 ( .A(n229), .B(n225), .C(n226), .D(n224), .S0(n245), .S1(
        Immediate_SE[9]), .Y(n126) );
  CLKINVX1 U219 ( .A(WBData[25]), .Y(n1049) );
  OA22X1 U220 ( .A0(n1072), .A1(n282), .B0(n1107), .B1(n279), .Y(n904) );
  NOR2XL U221 ( .A(n703), .B(n283), .Y(n105) );
  CLKINVX1 U222 ( .A(RData2[4]), .Y(n1105) );
  CLKINVX1 U223 ( .A(Immediate_SE[8]), .Y(n314) );
  CLKINVX1 U224 ( .A(n541), .Y(n982) );
  NAND2X1 U225 ( .A(n1020), .B(n328), .Y(n537) );
  NAND2X1 U226 ( .A(n1016), .B(n328), .Y(n992) );
  CLKINVX1 U227 ( .A(n383), .Y(n376) );
  MXI2X1 U228 ( .A(n184), .B(n182), .S0(Immediate_SE[7]), .Y(N501) );
  MXI2X1 U229 ( .A(n188), .B(n184), .S0(n309), .Y(N499) );
  AOI2BB1X1 U230 ( .A0N(n289), .A1N(n822), .B0(n821), .Y(n823) );
  MX2XL U231 ( .A(n397), .B(n396), .S0(n400), .Y(n406) );
  MX2XL U232 ( .A(n573), .B(n572), .S0(n581), .Y(n588) );
  NAND4X1 U233 ( .A(n124), .B(n877), .C(n876), .D(n875), .Y(next_ALUresult[5])
         );
  AOI22X1 U234 ( .A0(N337), .A1(n287), .B0(N209), .B1(n152), .Y(n124) );
  AOI22X1 U235 ( .A0(N345), .A1(n287), .B0(N217), .B1(n152), .Y(n119) );
  NAND4X1 U236 ( .A(n120), .B(n827), .C(n826), .D(n825), .Y(next_ALUresult[9])
         );
  AOI22X1 U237 ( .A0(N341), .A1(n287), .B0(N213), .B1(n152), .Y(n120) );
  MX2XL U238 ( .A(n963), .B(n962), .S0(n964), .Y(n971) );
  NOR2BX1 U239 ( .AN(n428), .B(n1013), .Y(n155) );
  INVX1 U240 ( .A(n310), .Y(n309) );
  CLKINVX1 U241 ( .A(n381), .Y(n940) );
  NAND3BX1 U242 ( .AN(n939), .B(n940), .C(n1013), .Y(n382) );
  CLKINVX1 U243 ( .A(n428), .Y(n380) );
  AOI211XL U244 ( .A0(Immediate_SE[2]), .A1(n443), .B0(ID_EX[3]), .C0(ID_EX[1]), .Y(n442) );
  NAND2XL U245 ( .A(Immediate_SE[5]), .B(n1119), .Y(n443) );
  INVX1 U246 ( .A(RData2[13]), .Y(n1096) );
  INVX1 U247 ( .A(RData2[15]), .Y(n1094) );
  INVX1 U248 ( .A(RData2[12]), .Y(n1097) );
  INVX1 U249 ( .A(RData2[8]), .Y(n1101) );
  INVX1 U250 ( .A(RData2[10]), .Y(n1099) );
  INVX1 U251 ( .A(RData2[9]), .Y(n1100) );
  INVX1 U252 ( .A(RData2[3]), .Y(n1106) );
  INVX1 U253 ( .A(RData2[5]), .Y(n1104) );
  INVX1 U254 ( .A(RData2[6]), .Y(n1103) );
  INVX1 U255 ( .A(RData2[7]), .Y(n1102) );
  NOR2XL U256 ( .A(n250), .B(n314), .Y(n107) );
  BUFX12 U257 ( .A(n935), .Y(n250) );
  MXI2X1 U258 ( .A(n241), .B(n8), .S0(Immediate_SE[8]), .Y(n165) );
  NAND2X1 U259 ( .A(n296), .B(n795), .Y(n792) );
  CLKINVX1 U260 ( .A(n329), .Y(n1110) );
  AO22X2 U261 ( .A0(N187), .A1(n148), .B0(N379), .B1(n150), .Y(n957) );
  MXI2X1 U262 ( .A(n178), .B(n169), .S0(Immediate_SE[7]), .Y(N505) );
  AO21X2 U263 ( .A0(N203), .A1(n1012), .B0(n154), .Y(n1022) );
  MXI2X1 U264 ( .A(n173), .B(n174), .S0(Immediate_SE[7]), .Y(N506) );
  NAND2XL U265 ( .A(ForwardA[1]), .B(n361), .Y(n931) );
  MXI2X1 U266 ( .A(n126), .B(n146), .S0(Immediate_SE[8]), .Y(n188) );
  MXI2X1 U267 ( .A(n202), .B(n194), .S0(Immediate_SE[7]), .Y(N495) );
  AOI2BB1X1 U268 ( .A0N(n290), .A1N(n909), .B0(n234), .Y(n910) );
  MXI2X1 U269 ( .A(n194), .B(n188), .S0(Immediate_SE[7]), .Y(N497) );
  AOI2BB1X1 U270 ( .A0N(n290), .A1N(n884), .B0(n235), .Y(n885) );
  AOI2BB1X1 U271 ( .A0N(n289), .A1N(n834), .B0(n833), .Y(n835) );
  MXI2X1 U272 ( .A(n199), .B(n191), .S0(Immediate_SE[7]), .Y(N496) );
  AOI2BB1X1 U273 ( .A0N(n290), .A1N(n897), .B0(n896), .Y(n898) );
  AOI2BB1X1 U274 ( .A0N(n289), .A1N(n847), .B0(n846), .Y(n848) );
  AOI2BB1X1 U275 ( .A0N(n289), .A1N(n859), .B0(n237), .Y(n860) );
  MXI2X1 U276 ( .A(n183), .B(n181), .S0(Immediate_SE[7]), .Y(N502) );
  AO22X1 U277 ( .A0(N172), .A1(n148), .B0(N364), .B1(n297), .Y(n946) );
  NAND2X1 U278 ( .A(n149), .B(n954), .Y(n951) );
  NAND2X1 U279 ( .A(n296), .B(n755), .Y(n752) );
  MX2XL U280 ( .A(n498), .B(n496), .S0(n507), .Y(n517) );
  MX2XL U281 ( .A(n436), .B(n432), .S0(n449), .Y(n462) );
  MX2XL U282 ( .A(n413), .B(n412), .S0(n416), .Y(n423) );
  MX2XL U283 ( .A(n994), .B(n993), .S0(n996), .Y(n1005) );
  MX2XL U284 ( .A(n471), .B(n469), .S0(n478), .Y(n489) );
  MX2XL U285 ( .A(n526), .B(n525), .S0(n534), .Y(n548) );
  MX2XL U286 ( .A(n556), .B(n555), .S0(n561), .Y(n567) );
  MX2XL U287 ( .A(n375), .B(n374), .S0(n385), .Y(n391) );
  NAND2XL U288 ( .A(ForwardA[0]), .B(n362), .Y(n930) );
  CLKMX2X2 U289 ( .A(n189), .B(n8), .S0(n245), .Y(n125) );
  INVXL U290 ( .A(n252), .Y(n998) );
  INVX1 U291 ( .A(WBData[28]), .Y(n1046) );
  INVX1 U292 ( .A(WBData[29]), .Y(n1045) );
  NAND3BXL U293 ( .AN(n380), .B(n940), .C(n1013), .Y(n1009) );
  INVX3 U294 ( .A(n318), .Y(n317) );
  NAND3BXL U295 ( .AN(n1014), .B(n381), .C(n1013), .Y(n379) );
  NAND3BXL U296 ( .AN(n1014), .B(n155), .C(n381), .Y(n373) );
  AND2XL U297 ( .A(n381), .B(n380), .Y(n159) );
  AND2XL U298 ( .A(n153), .B(n381), .Y(n160) );
  AND2XL U299 ( .A(n1013), .B(n380), .Y(n161) );
  NAND2X1 U300 ( .A(RData1[1]), .B(n6), .Y(n915) );
  NAND2X1 U301 ( .A(RData1[4]), .B(n6), .Y(n878) );
  NAND2XL U302 ( .A(RData1[3]), .B(n6), .Y(n890) );
  MX2XL U303 ( .A(n1011), .B(n1010), .S0(n1015), .Y(n1024) );
  CLKINVX1 U304 ( .A(RData2[2]), .Y(n1107) );
  CLKINVX1 U305 ( .A(RData2[1]), .Y(n1040) );
  CLKINVX1 U306 ( .A(RData2[0]), .Y(n1036) );
  AND2XL U307 ( .A(n185), .B(n980), .Y(n456) );
  AND2XL U308 ( .A(n168), .B(n980), .Y(n419) );
  AO22X2 U309 ( .A0(N198), .A1(n298), .B0(N390), .B1(n297), .Y(n403) );
  MXI2XL U310 ( .A(n244), .B(n144), .S0(Immediate_SE[8]), .Y(n194) );
  INVXL U311 ( .A(n230), .Y(n244) );
  AOI2BB1XL U312 ( .A0N(n139), .A1N(n995), .B0(n109), .Y(n1003) );
  INVXL U313 ( .A(n313), .Y(n729) );
  AOI2BB1XL U314 ( .A0N(n1020), .A1N(n1019), .B0(n1018), .Y(n1021) );
  AO22X2 U315 ( .A0(N195), .A1(n298), .B0(N387), .B1(n297), .Y(n484) );
  INVXL U316 ( .A(n214), .Y(n513) );
  INVXL U317 ( .A(n231), .Y(n544) );
  MXI3XL U318 ( .A(n164), .B(n165), .C(n1018), .S0(Immediate_SE[7]), .S1(
        Immediate_SE[10]), .Y(N508) );
  AOI2BB1XL U319 ( .A0N(n289), .A1N(n809), .B0(n808), .Y(n810) );
  AO22X2 U320 ( .A0(N191), .A1(n298), .B0(N383), .B1(n297), .Y(n585) );
  AOI2BB1XL U321 ( .A0N(n290), .A1N(n872), .B0(n236), .Y(n873) );
  AOI2BB2XL U322 ( .B0(n285), .B1(n378), .A0N(n995), .A1N(n377), .Y(n389) );
  INVXL U323 ( .A(n140), .Y(n377) );
  AOI2BB1XL U324 ( .A0N(n1000), .A1N(n979), .B0(n256), .Y(n984) );
  AOI2BB1XL U325 ( .A0N(n1000), .A1N(n966), .B0(n258), .Y(n967) );
  OA22XL U326 ( .A0(n198), .A1(n257), .B0(n186), .B1(n256), .Y(n477) );
  OA22XL U327 ( .A0(n158), .A1(n727), .B0(n130), .B1(n725), .Y(n474) );
  OA22XL U328 ( .A0(n220), .A1(n258), .B0(n157), .B1(n728), .Y(n475) );
  OA22XL U329 ( .A0(n139), .A1(n724), .B0(n177), .B1(n621), .Y(n472) );
  OA22XL U330 ( .A0(n256), .A1(n248), .B0(n232), .B1(n258), .Y(n576) );
  NOR2X1 U331 ( .A(n311), .B(n309), .Y(n353) );
  NAND2X1 U332 ( .A(n349), .B(n353), .Y(n215) );
  NAND2X1 U333 ( .A(n350), .B(n353), .Y(n232) );
  AOI2BB1XL U334 ( .A0N(n290), .A1N(n450), .B0(n724), .Y(n452) );
  AOI2BB1XL U335 ( .A0N(n1000), .A1N(n417), .B0(n725), .Y(n418) );
  AOI2BB1XL U336 ( .A0N(n1000), .A1N(n386), .B0(n728), .Y(n387) );
  NAND2XL U337 ( .A(n149), .B(n256), .Y(n975) );
  NAND2XL U338 ( .A(n296), .B(n258), .Y(n962) );
  NAND2XL U339 ( .A(n296), .B(n781), .Y(n778) );
  NAND2XL U340 ( .A(n296), .B(n728), .Y(n374) );
  NAND2XL U341 ( .A(n296), .B(n621), .Y(n469) );
  NAND2XL U342 ( .A(n296), .B(n724), .Y(n432) );
  NAND2XL U343 ( .A(n296), .B(n768), .Y(n765) );
  NAND2XL U344 ( .A(n296), .B(n725), .Y(n412) );
  NAND2XL U345 ( .A(n161), .B(n1018), .Y(n1010) );
  NAND2X1 U346 ( .A(n348), .B(n358), .Y(n198) );
  NAND2X1 U347 ( .A(n351), .B(n359), .Y(n157) );
  NAND2X1 U348 ( .A(n354), .B(n358), .Y(n158) );
  NOR3BX1 U349 ( .AN(n1003), .B(n1002), .C(n1001), .Y(n1004) );
  NOR3BX1 U350 ( .AN(n389), .B(n388), .C(n387), .Y(n390) );
  AOI22X1 U351 ( .A0(N347), .A1(n287), .B0(N219), .B1(n286), .Y(n110) );
  AOI22X1 U352 ( .A0(N346), .A1(n287), .B0(N218), .B1(n286), .Y(n111) );
  AOI22X1 U353 ( .A0(N343), .A1(n287), .B0(N215), .B1(n286), .Y(n112) );
  AOI22X1 U354 ( .A0(N332), .A1(n287), .B0(N204), .B1(n152), .Y(n113) );
  AOI22X1 U355 ( .A0(N342), .A1(n287), .B0(N214), .B1(n286), .Y(n114) );
  AOI22X1 U356 ( .A0(N344), .A1(n287), .B0(N216), .B1(n152), .Y(n115) );
  AOI22X1 U357 ( .A0(N339), .A1(n287), .B0(N211), .B1(n152), .Y(n116) );
  AOI22X1 U358 ( .A0(N340), .A1(n287), .B0(N212), .B1(n152), .Y(n117) );
  AOI22X1 U359 ( .A0(N338), .A1(n287), .B0(N210), .B1(n152), .Y(n118) );
  INVXL U360 ( .A(n156), .Y(n398) );
  MXI2XL U361 ( .A(ALUData2[15]), .B(n271), .S0(n307), .Y(n216) );
  MXI2XL U362 ( .A(n262), .B(n261), .S0(Immediate_SE[6]), .Y(n213) );
  MXI2XL U363 ( .A(n271), .B(n270), .S0(Immediate_SE[6]), .Y(n221) );
  MXI2XL U364 ( .A(n270), .B(n267), .S0(Immediate_SE[6]), .Y(n210) );
  MXI2XL U365 ( .A(n264), .B(n263), .S0(Immediate_SE[6]), .Y(n208) );
  MXI2XL U366 ( .A(n265), .B(n264), .S0(n249), .Y(n218) );
  MXI2XL U367 ( .A(n266), .B(n265), .S0(Immediate_SE[6]), .Y(n212) );
  MXI2XL U368 ( .A(ALUData2[8]), .B(ALUData2[9]), .S0(n249), .Y(n227) );
  MXI2XL U369 ( .A(n267), .B(n266), .S0(n249), .Y(n223) );
  MXI2XL U370 ( .A(n260), .B(n259), .S0(Immediate_SE[6]), .Y(n209) );
  MXI2XL U371 ( .A(n261), .B(n260), .S0(Immediate_SE[6]), .Y(n219) );
  MXI2XL U372 ( .A(n253), .B(n252), .S0(Immediate_SE[6]), .Y(n207) );
  MXI2XL U373 ( .A(n254), .B(n253), .S0(n307), .Y(n217) );
  MXI2XL U374 ( .A(n255), .B(n254), .S0(Immediate_SE[6]), .Y(n211) );
  MXI2XL U375 ( .A(n259), .B(n255), .S0(n249), .Y(n222) );
  MXI2XL U376 ( .A(n263), .B(n262), .S0(n249), .Y(n225) );
  MXI2XL U377 ( .A(n252), .B(n251), .S0(n249), .Y(n224) );
  INVX1 U378 ( .A(n259), .Y(n727) );
  INVX1 U379 ( .A(n263), .Y(n620) );
  INVX1 U380 ( .A(n264), .Y(n624) );
  AOI22X1 U381 ( .A0(N335), .A1(n287), .B0(N207), .B1(n152), .Y(n121) );
  AOI22X1 U382 ( .A0(N334), .A1(n151), .B0(N206), .B1(n286), .Y(n122) );
  INVX1 U383 ( .A(n265), .Y(n623) );
  MXI2XL U384 ( .A(n243), .B(n251), .S0(n245), .Y(n174) );
  INVXL U385 ( .A(n266), .Y(n582) );
  AO22XL U386 ( .A0(n259), .A1(n981), .B0(n255), .B1(n499), .Y(n415) );
  MXI4X1 U387 ( .A(n228), .B(n213), .C(n216), .D(n1018), .S0(n245), .S1(n246), 
        .Y(n127) );
  MXI3XL U388 ( .A(n240), .B(n10), .C(n251), .S0(Immediate_SE[8]), .S1(n245), 
        .Y(n170) );
  INVX1 U389 ( .A(n176), .Y(n240) );
  AO22XL U390 ( .A0(n259), .A1(n731), .B0(n255), .B1(n730), .Y(n502) );
  AO22XL U391 ( .A0(n259), .A1(n730), .B0(n255), .B1(n1115), .Y(n529) );
  AO22XL U392 ( .A0(n261), .A1(n499), .B0(n260), .B1(n1111), .Y(n504) );
  MXI3XL U393 ( .A(n921), .B(n234), .C(n204), .S0(n249), .S1(n315), .Y(n203)
         );
  AO22XL U394 ( .A0(n1115), .A1(n263), .B0(n1112), .B1(n262), .Y(n732) );
  AO22XL U395 ( .A0(n271), .A1(n1114), .B0(n270), .B1(n981), .Y(n735) );
  AND2XL U396 ( .A(n376), .B(n251), .Y(n154) );
  NOR3X1 U397 ( .A(n317), .B(n307), .C(n316), .Y(n349) );
  NOR3X1 U398 ( .A(n316), .B(n317), .C(n308), .Y(n350) );
  NOR2X1 U399 ( .A(n310), .B(n314), .Y(n348) );
  NOR2X1 U400 ( .A(n310), .B(n311), .Y(n354) );
  NOR2X1 U401 ( .A(n314), .B(n309), .Y(n351) );
  INVXL U402 ( .A(ALUData1[22]), .Y(n507) );
  INVXL U403 ( .A(ALUData1[23]), .Y(n478) );
  INVXL U404 ( .A(ALUData1[27]), .Y(n385) );
  INVXL U405 ( .A(ALUData1[29]), .Y(n977) );
  INVXL U406 ( .A(ALUData1[26]), .Y(n400) );
  INVXL U407 ( .A(ALUData1[30]), .Y(n996) );
  INVXL U408 ( .A(ALUData1[31]), .Y(n1015) );
  INVXL U409 ( .A(ALUData1[16]), .Y(n737) );
  INVXL U410 ( .A(ALUData1[28]), .Y(n964) );
  INVXL U411 ( .A(ALUData1[0]), .Y(n942) );
  AOI2BB1XL U412 ( .A0N(n262), .A1N(n294), .B0(n289), .Y(n471) );
  AOI2BB1XL U413 ( .A0N(n263), .A1N(n294), .B0(n289), .Y(n498) );
  AOI2BB1XL U414 ( .A0N(n261), .A1N(n291), .B0(n289), .Y(n436) );
  AOI2BB1XL U415 ( .A0N(n264), .A1N(n294), .B0(n289), .Y(n526) );
  AOI2BB1XL U416 ( .A0N(n260), .A1N(n291), .B0(n289), .Y(n413) );
  AOI2BB1XL U417 ( .A0N(n271), .A1N(n291), .B0(n288), .Y(n723) );
  AOI2BB1XL U418 ( .A0N(n259), .A1N(n294), .B0(n288), .Y(n397) );
  AOI2BB1XL U419 ( .A0N(n265), .A1N(n294), .B0(n288), .Y(n556) );
  AOI2BB1XL U420 ( .A0N(n267), .A1N(n294), .B0(n288), .Y(n594) );
  AOI2BB1XL U421 ( .A0N(n266), .A1N(n294), .B0(n288), .Y(n573) );
  AOI2BB1XL U422 ( .A0N(n252), .A1N(n291), .B0(n288), .Y(n994) );
  AOI2BB1XL U423 ( .A0N(n270), .A1N(n294), .B0(n288), .Y(n619) );
  AOI2BB1XL U424 ( .A0N(n255), .A1N(n291), .B0(n288), .Y(n375) );
  AOI2BB1XL U425 ( .A0N(n254), .A1N(n992), .B0(n288), .Y(n963) );
  AOI2BB1XL U426 ( .A0N(n253), .A1N(n291), .B0(n290), .Y(n976) );
  INVXL U427 ( .A(n271), .Y(n738) );
  AOI2BB1XL U428 ( .A0N(n251), .A1N(n1009), .B0(n1020), .Y(n1011) );
  INVXL U429 ( .A(n267), .Y(n606) );
  INVXL U430 ( .A(n270), .Y(n677) );
  INVX1 U431 ( .A(n314), .Y(n311) );
  AO22XL U432 ( .A0(n313), .A1(n252), .B0(n312), .B1(n251), .Y(n627) );
  AND3XL U433 ( .A(n285), .B(n252), .C(n981), .Y(n983) );
  INVX1 U434 ( .A(n316), .Y(n315) );
  NAND2X1 U435 ( .A(n549), .B(n328), .Y(n451) );
  NAND2BX1 U436 ( .AN(ForwardB[0]), .B(n347), .Y(n355) );
  AOI2BB2XL U437 ( .B0(Immediate_SE[15]), .B1(n789), .A0N(n1156), .A1N(n283), 
        .Y(n748) );
  OA22XL U438 ( .A0(n1068), .A1(n282), .B0(n1103), .B1(n279), .Y(n854) );
  AOI2BB2XL U439 ( .B0(Immediate_SE[14]), .B1(n789), .A0N(n1168), .A1N(n283), 
        .Y(n750) );
  OA22XL U440 ( .A0(n1067), .A1(n282), .B0(n1102), .B1(n279), .Y(n841) );
  NAND2XL U441 ( .A(RData1[18]), .B(n6), .Y(n591) );
  NAND2XL U442 ( .A(RData1[23]), .B(n6), .Y(n466) );
  NAND2XL U443 ( .A(RData1[19]), .B(n6), .Y(n570) );
  NAND2XL U444 ( .A(RData1[21]), .B(n6), .Y(n522) );
  NAND2XL U445 ( .A(RData1[17]), .B(n6), .Y(n615) );
  NAND2XL U446 ( .A(RData1[14]), .B(n6), .Y(n749) );
  NAND2XL U447 ( .A(RData1[26]), .B(n6), .Y(n394) );
  NAND2XL U448 ( .A(RData1[13]), .B(n6), .Y(n762) );
  NAND2XL U449 ( .A(RData1[15]), .B(n6), .Y(n747) );
  NAND2XL U450 ( .A(RData1[5]), .B(n6), .Y(n865) );
  NAND2XL U451 ( .A(RData1[8]), .B(n6), .Y(n828) );
  NAND2XL U452 ( .A(RData1[16]), .B(n6), .Y(n719) );
  NAND2XL U453 ( .A(RData1[12]), .B(n6), .Y(n775) );
  NAND2XL U454 ( .A(RData1[2]), .B(n6), .Y(n903) );
  NAND2XL U455 ( .A(RData1[27]), .B(n6), .Y(n370) );
  NAND2XL U456 ( .A(RData1[29]), .B(n6), .Y(n366) );
  NAND2XL U457 ( .A(RData1[30]), .B(n6), .Y(n365) );
  NAND2XL U458 ( .A(RData1[31]), .B(n6), .Y(n363) );
  NAND2XL U459 ( .A(RData1[28]), .B(n6), .Y(n369) );
  AOI211XL U460 ( .A0(Immediate_SE[1]), .A1(n1118), .B0(Immediate_SE[4]), .C0(
        ID_EX[1]), .Y(n445) );
  NAND3XL U461 ( .A(Immediate_SE[5]), .B(n439), .C(n445), .Y(n444) );
  AOI2BB1XL U462 ( .A0N(Immediate_SE[2]), .A1N(n1120), .B0(Immediate_SE[3]), 
        .Y(n439) );
  OAI211XL U463 ( .A0(Immediate_SE[5]), .A1(n431), .B0(n1116), .C0(n433), .Y(
        n429) );
  AOI211XL U464 ( .A0(Immediate_SE[1]), .A1(n1120), .B0(Immediate_SE[3]), .C0(
        Immediate_SE[2]), .Y(n431) );
  INVXL U465 ( .A(Immediate_SE[3]), .Y(n1117) );
  INVXL U466 ( .A(Immediate_SE[4]), .Y(n1116) );
  INVX1 U467 ( .A(RData2[14]), .Y(n1095) );
  INVX1 U468 ( .A(RData2[16]), .Y(n1093) );
  AO21XL U469 ( .A0(Immediate_SE[0]), .A1(Immediate_SE[5]), .B0(n1119), .Y(
        n435) );
  OA22XL U470 ( .A0(n302), .A1(n710), .B0(n333), .B1(n1037), .Y(n1038) );
  OAI2BB1XL U471 ( .A0N(RegisterRd[1]), .A1N(n321), .B0(n128), .Y(n1076) );
  AOI22XL U472 ( .A0(ID_RegisterRt[1]), .A1(n162), .B0(ID_RegisterRd[1]), .B1(
        n163), .Y(n128) );
  OAI2BB1XL U473 ( .A0N(n322), .A1N(RegisterRd[4]), .B0(n131), .Y(n1073) );
  AOI22XL U474 ( .A0(ID_RegisterRt[4]), .A1(n162), .B0(ID_RegisterRd[4]), .B1(
        n163), .Y(n131) );
  AO21XL U475 ( .A0(RegisterRd[3]), .A1(n322), .B0(n1032), .Y(n1074) );
  AO22XL U476 ( .A0(ID_RegisterRt[3]), .A1(n162), .B0(ID_RegisterRd[3]), .B1(
        n163), .Y(n1032) );
  OAI2BB1XL U477 ( .A0N(n322), .A1N(RegisterRd[0]), .B0(n132), .Y(n1077) );
  AOI22XL U478 ( .A0(ID_RegisterRt[0]), .A1(n162), .B0(ID_RegisterRd[0]), .B1(
        n163), .Y(n132) );
  OAI2BB1XL U479 ( .A0N(n322), .A1N(RegisterRd[2]), .B0(n133), .Y(n1075) );
  AOI22XL U480 ( .A0(ID_RegisterRt[2]), .A1(n162), .B0(ID_RegisterRd[2]), .B1(
        n163), .Y(n133) );
  XNOR2XL U481 ( .A(ForwardB[0]), .B(ForwardB[1]), .Y(n549) );
  NAND3BXL U482 ( .AN(ForwardB[1]), .B(n328), .C(ForwardB[0]), .Y(n453) );
  NAND3BXL U483 ( .AN(ForwardB[0]), .B(ForwardB[1]), .C(n328), .Y(n455) );
  OAI221X4 U484 ( .A0(n1063), .A1(n281), .B0(n1098), .B1(n280), .C0(n790), .Y(
        n134) );
  AOI2BB2XL U485 ( .B0(Immediate_SE[11]), .B1(n789), .A0N(n1165), .A1N(n283), 
        .Y(n790) );
  CLKBUFX3 U486 ( .A(n982), .Y(n284) );
  CLKBUFX3 U487 ( .A(n982), .Y(n285) );
  CLKBUFX3 U488 ( .A(n991), .Y(n288) );
  CLKBUFX3 U489 ( .A(n991), .Y(n289) );
  CLKBUFX3 U490 ( .A(n991), .Y(n290) );
  INVX3 U491 ( .A(n291), .Y(n293) );
  INVX3 U492 ( .A(n291), .Y(n292) );
  CLKBUFX3 U493 ( .A(n291), .Y(n294) );
  CLKBUFX3 U494 ( .A(n933), .Y(n282) );
  CLKBUFX3 U495 ( .A(n932), .Y(n278) );
  NAND2X1 U496 ( .A(n376), .B(n324), .Y(n541) );
  CLKINVX1 U497 ( .A(n537), .Y(n991) );
  NOR2X1 U498 ( .A(n140), .B(n1111), .Y(n129) );
  NOR2X1 U499 ( .A(n295), .B(n1110), .Y(n268) );
  NOR2X1 U500 ( .A(n168), .B(n730), .Y(n156) );
  CLKBUFX3 U501 ( .A(n992), .Y(n291) );
  CLKINVX1 U502 ( .A(n323), .Y(n322) );
  CLKINVX1 U503 ( .A(n731), .Y(n597) );
  CLKINVX1 U504 ( .A(n1111), .Y(n622) );
  CLKINVX1 U505 ( .A(n177), .Y(n1114) );
  CLKINVX1 U506 ( .A(n1115), .Y(n596) );
  INVX3 U507 ( .A(n324), .Y(n321) );
  INVX3 U508 ( .A(n325), .Y(n320) );
  CLKINVX1 U509 ( .A(n1112), .Y(n575) );
  CLKINVX1 U510 ( .A(n625), .Y(n574) );
  CLKINVX1 U511 ( .A(n295), .Y(n595) );
  INVX3 U512 ( .A(n326), .Y(n319) );
  MXI2X1 U513 ( .A(n147), .B(n136), .S0(Immediate_SE[8]), .Y(n183) );
  MXI2X1 U514 ( .A(n239), .B(n9), .S0(n311), .Y(n164) );
  CLKINVX1 U515 ( .A(n180), .Y(n239) );
  AO22X1 U516 ( .A0(N356), .A1(n151), .B0(N228), .B1(n286), .Y(n465) );
  AO22X1 U517 ( .A0(N357), .A1(n151), .B0(N229), .B1(n286), .Y(n425) );
  AO22X1 U518 ( .A0(N358), .A1(n151), .B0(N230), .B1(n286), .Y(n408) );
  AO22X1 U519 ( .A0(N359), .A1(n151), .B0(N231), .B1(n286), .Y(n393) );
  AO22X1 U520 ( .A0(N353), .A1(n151), .B0(N225), .B1(n286), .Y(n551) );
  AO22X1 U521 ( .A0(N355), .A1(n151), .B0(N227), .B1(n286), .Y(n492) );
  AO22X1 U522 ( .A0(N352), .A1(n151), .B0(N224), .B1(n286), .Y(n569) );
  AO22X1 U523 ( .A0(N351), .A1(n287), .B0(N223), .B1(n286), .Y(n590) );
  AO22X1 U524 ( .A0(N354), .A1(n151), .B0(N226), .B1(n286), .Y(n520) );
  AO22X1 U525 ( .A0(N350), .A1(n287), .B0(N222), .B1(n286), .Y(n614) );
  CLKBUFX3 U526 ( .A(n931), .Y(n275) );
  CLKBUFX3 U527 ( .A(n931), .Y(n276) );
  MXI2X1 U528 ( .A(n146), .B(n145), .S0(Immediate_SE[8]), .Y(n182) );
  NAND2X1 U529 ( .A(n129), .B(n130), .Y(n106) );
  CLKINVX1 U530 ( .A(n172), .Y(n241) );
  NAND2BX1 U531 ( .AN(n185), .B(n186), .Y(n168) );
  NAND2X1 U532 ( .A(n156), .B(n157), .Y(n140) );
  NAND2BX1 U533 ( .AN(n231), .B(n232), .Y(n214) );
  NAND2BX1 U534 ( .AN(n214), .B(n215), .Y(n197) );
  NAND2BX1 U535 ( .AN(n197), .B(n198), .Y(n185) );
  NAND2BX1 U536 ( .AN(n247), .B(n248), .Y(n231) );
  NAND2X1 U537 ( .A(n330), .B(n331), .Y(n312) );
  NAND2X1 U538 ( .A(n268), .B(n269), .Y(n247) );
  CLKBUFX3 U539 ( .A(n335), .Y(n326) );
  CLKBUFX3 U540 ( .A(n335), .Y(n327) );
  CLKBUFX3 U541 ( .A(n335), .Y(n325) );
  CLKBUFX3 U542 ( .A(n336), .Y(n323) );
  CLKBUFX3 U543 ( .A(n336), .Y(n324) );
  CLKBUFX3 U544 ( .A(n334), .Y(n328) );
  CLKBUFX3 U545 ( .A(n334), .Y(n332) );
  CLKBUFX3 U546 ( .A(n148), .Y(n298) );
  CLKBUFX3 U547 ( .A(n150), .Y(n297) );
  CLKBUFX3 U548 ( .A(n997), .Y(n299) );
  CLKBUFX3 U549 ( .A(n997), .Y(n300) );
  CLKBUFX3 U550 ( .A(n149), .Y(n296) );
  CLKBUFX3 U551 ( .A(n151), .Y(n287) );
  CLKBUFX3 U552 ( .A(n152), .Y(n286) );
  NAND2X1 U553 ( .A(n359), .B(n353), .Y(n177) );
  CLKINVX1 U554 ( .A(n130), .Y(n1113) );
  CLKINVX1 U555 ( .A(n157), .Y(n731) );
  CLKINVX1 U556 ( .A(n220), .Y(n730) );
  CLKINVX1 U557 ( .A(n130), .Y(n499) );
  CLKINVX1 U558 ( .A(n158), .Y(n1111) );
  CLKINVX1 U559 ( .A(n232), .Y(n626) );
  CLKINVX1 U560 ( .A(n215), .Y(n625) );
  CLKINVX1 U561 ( .A(n198), .Y(n1112) );
  CLKINVX1 U562 ( .A(n186), .Y(n1115) );
  INVX3 U563 ( .A(n139), .Y(n981) );
  CLKBUFX3 U564 ( .A(n317), .Y(n245) );
  CLKBUFX3 U565 ( .A(n315), .Y(n246) );
  CLKBUFX3 U566 ( .A(n307), .Y(n249) );
  CLKBUFX3 U567 ( .A(n334), .Y(n333) );
  CLKINVX1 U568 ( .A(n248), .Y(n1109) );
  CLKINVX1 U569 ( .A(n269), .Y(n1108) );
  CLKBUFX3 U570 ( .A(n339), .Y(n341) );
  CLKBUFX3 U571 ( .A(n339), .Y(n342) );
  CLKBUFX3 U572 ( .A(n338), .Y(n343) );
  CLKBUFX3 U573 ( .A(n338), .Y(n344) );
  CLKBUFX3 U574 ( .A(n338), .Y(n345) );
  CLKBUFX3 U575 ( .A(n339), .Y(n346) );
  NAND2X1 U576 ( .A(n352), .B(n355), .Y(n933) );
  CLKINVX1 U577 ( .A(n355), .Y(n357) );
  CLKINVX1 U578 ( .A(n356), .Y(n352) );
  NAND2X1 U579 ( .A(n356), .B(n355), .Y(n935) );
  AOI211X1 U580 ( .A0(N508), .A1(n284), .B0(n957), .C0(n956), .Y(n958) );
  AOI2BB1X1 U581 ( .A0N(n290), .A1N(n955), .B0(n954), .Y(n956) );
  AOI211X1 U582 ( .A0(N507), .A1(n285), .B0(n758), .C0(n757), .Y(n759) );
  AOI2BB1X1 U583 ( .A0N(n289), .A1N(n756), .B0(n755), .Y(n757) );
  MXI2X1 U584 ( .A(n169), .B(n170), .S0(Immediate_SE[7]), .Y(N507) );
  AO22X1 U585 ( .A0(N186), .A1(n298), .B0(N378), .B1(n297), .Y(n758) );
  AOI211X1 U586 ( .A0(N506), .A1(n285), .B0(n771), .C0(n770), .Y(n772) );
  AOI2BB1X1 U587 ( .A0N(n289), .A1N(n769), .B0(n768), .Y(n770) );
  AOI211X1 U588 ( .A0(N505), .A1(n285), .B0(n784), .C0(n783), .Y(n785) );
  AOI2BB1X1 U589 ( .A0N(n289), .A1N(n782), .B0(n781), .Y(n783) );
  AO22X1 U590 ( .A0(N184), .A1(n298), .B0(N376), .B1(n297), .Y(n784) );
  AOI211X1 U591 ( .A0(N504), .A1(n285), .B0(n798), .C0(n797), .Y(n799) );
  AOI2BB1X1 U592 ( .A0N(n289), .A1N(n796), .B0(n795), .Y(n797) );
  MXI2X1 U593 ( .A(n181), .B(n173), .S0(Immediate_SE[7]), .Y(N504) );
  AO22X1 U594 ( .A0(N183), .A1(n298), .B0(N375), .B1(n297), .Y(n798) );
  AOI211X1 U595 ( .A0(N503), .A1(n285), .B0(n811), .C0(n810), .Y(n812) );
  MXI2X1 U596 ( .A(n182), .B(n178), .S0(Immediate_SE[7]), .Y(N503) );
  AO22X1 U597 ( .A0(N182), .A1(n298), .B0(N374), .B1(n297), .Y(n811) );
  AOI211X1 U598 ( .A0(N502), .A1(n285), .B0(n824), .C0(n823), .Y(n825) );
  AO22X1 U599 ( .A0(N181), .A1(n298), .B0(N373), .B1(n297), .Y(n824) );
  AOI211X1 U600 ( .A0(N501), .A1(n285), .B0(n836), .C0(n835), .Y(n837) );
  AO22X1 U601 ( .A0(N180), .A1(n298), .B0(N372), .B1(n150), .Y(n836) );
  AOI211X1 U602 ( .A0(N500), .A1(n285), .B0(n849), .C0(n848), .Y(n850) );
  MXI2X1 U603 ( .A(n187), .B(n183), .S0(Immediate_SE[7]), .Y(N500) );
  AOI211X1 U604 ( .A0(N499), .A1(n285), .B0(n861), .C0(n860), .Y(n862) );
  AO22X1 U605 ( .A0(N178), .A1(n148), .B0(N370), .B1(n150), .Y(n861) );
  AOI211X1 U606 ( .A0(N498), .A1(n285), .B0(n874), .C0(n873), .Y(n875) );
  AO22X1 U607 ( .A0(N177), .A1(n148), .B0(N369), .B1(n297), .Y(n874) );
  AOI211X1 U608 ( .A0(N495), .A1(n284), .B0(n911), .C0(n910), .Y(n912) );
  AO22X1 U609 ( .A0(N174), .A1(n148), .B0(N366), .B1(n150), .Y(n911) );
  AOI211X1 U610 ( .A0(N494), .A1(n284), .B0(n924), .C0(n923), .Y(n925) );
  AOI2BB1X1 U611 ( .A0N(n290), .A1N(n922), .B0(n921), .Y(n923) );
  MXI2X1 U612 ( .A(n205), .B(n199), .S0(Immediate_SE[7]), .Y(N494) );
  AO22X1 U613 ( .A0(N173), .A1(n148), .B0(N365), .B1(n150), .Y(n924) );
  AOI211X1 U614 ( .A0(N497), .A1(n284), .B0(n886), .C0(n885), .Y(n887) );
  AO22X1 U615 ( .A0(N176), .A1(n148), .B0(N368), .B1(n150), .Y(n886) );
  AOI211X1 U616 ( .A0(N496), .A1(n285), .B0(n899), .C0(n898), .Y(n900) );
  AO22X1 U617 ( .A0(N175), .A1(n148), .B0(N367), .B1(n150), .Y(n899) );
  CLKMX2X2 U618 ( .A(n216), .B(n213), .S0(n246), .Y(n180) );
  AOI211X1 U619 ( .A0(N395), .A1(n159), .B0(n1022), .C0(n1021), .Y(n1023) );
  MXI2X1 U620 ( .A(n137), .B(n175), .S0(Immediate_SE[8]), .Y(n178) );
  MXI2X1 U621 ( .A(n176), .B(n1018), .S0(n245), .Y(n175) );
  MXI2X1 U622 ( .A(n138), .B(n179), .S0(Immediate_SE[8]), .Y(n181) );
  MXI2X1 U623 ( .A(n180), .B(n1018), .S0(n317), .Y(n179) );
  MXI2X1 U624 ( .A(n136), .B(n171), .S0(Immediate_SE[8]), .Y(n173) );
  MXI2X1 U625 ( .A(n172), .B(n1018), .S0(n245), .Y(n171) );
  MXI2X1 U626 ( .A(n127), .B(n138), .S0(Immediate_SE[8]), .Y(n187) );
  MXI2X1 U627 ( .A(n125), .B(n147), .S0(Immediate_SE[8]), .Y(n191) );
  MXI2X1 U628 ( .A(n192), .B(n10), .S0(n245), .Y(n230) );
  MXI3X1 U629 ( .A(n195), .B(n9), .C(n127), .S0(n245), .S1(Immediate_SE[8]), 
        .Y(n199) );
  MXI3X1 U630 ( .A(n896), .B(n235), .C(n196), .S0(n249), .S1(n246), .Y(n195)
         );
  MXI3X1 U631 ( .A(n200), .B(n242), .C(n126), .S0(Immediate_SE[10]), .S1(
        Immediate_SE[8]), .Y(n202) );
  CLKINVX1 U632 ( .A(n167), .Y(n242) );
  MXI3X1 U633 ( .A(n234), .B(n896), .C(n201), .S0(n249), .S1(Immediate_SE[9]), 
        .Y(n200) );
  MXI4X1 U634 ( .A(n190), .B(n207), .C(n208), .D(n1018), .S0(n245), .S1(n246), 
        .Y(n136) );
  MXI4X1 U635 ( .A(n193), .B(n217), .C(n218), .D(n1018), .S0(n245), .S1(n246), 
        .Y(n137) );
  MXI4X1 U636 ( .A(n196), .B(n211), .C(n212), .D(n1018), .S0(n245), .S1(n246), 
        .Y(n138) );
  AO22X1 U637 ( .A0(N199), .A1(n148), .B0(N391), .B1(n150), .Y(n388) );
  AO22X1 U638 ( .A0(N202), .A1(n298), .B0(N394), .B1(n297), .Y(n1002) );
  AO22X1 U639 ( .A0(N190), .A1(n298), .B0(N382), .B1(n297), .Y(n609) );
  AO22X1 U640 ( .A0(N188), .A1(n298), .B0(N380), .B1(n297), .Y(n741) );
  AO22X1 U641 ( .A0(N192), .A1(n298), .B0(N384), .B1(n297), .Y(n564) );
  AO22X1 U642 ( .A0(N189), .A1(n298), .B0(N381), .B1(n297), .Y(n713) );
  AO22X1 U643 ( .A0(N200), .A1(n148), .B0(N392), .B1(n150), .Y(n968) );
  AO22X1 U644 ( .A0(N196), .A1(n298), .B0(N388), .B1(n297), .Y(n459) );
  AO22X1 U645 ( .A0(N201), .A1(n148), .B0(N393), .B1(n150), .Y(n985) );
  AO22X1 U646 ( .A0(N197), .A1(n298), .B0(N389), .B1(n297), .Y(n421) );
  AO22X1 U647 ( .A0(N362), .A1(n287), .B0(N234), .B1(n152), .Y(n1007) );
  AO22X1 U648 ( .A0(N360), .A1(n151), .B0(N232), .B1(n286), .Y(n973) );
  AO22X1 U649 ( .A0(N361), .A1(n151), .B0(N233), .B1(n286), .Y(n989) );
  AO22X1 U650 ( .A0(N363), .A1(n160), .B0(N235), .B1(n1008), .Y(n1025) );
  AO22X1 U651 ( .A0(N348), .A1(n287), .B0(N220), .B1(n286), .Y(n746) );
  AO22X1 U652 ( .A0(N349), .A1(n151), .B0(N221), .B1(n286), .Y(n718) );
  CLKBUFX3 U653 ( .A(n272), .Y(n274) );
  CLKBUFX3 U654 ( .A(n930), .Y(n272) );
  NAND2X1 U655 ( .A(n154), .B(n323), .Y(n995) );
  OAI222XL U656 ( .A0(n215), .A1(n256), .B0(n232), .B1(n257), .C0(n198), .C1(
        n258), .Y(n528) );
  OAI222XL U657 ( .A0(n198), .A1(n256), .B0(n215), .B1(n257), .C0(n186), .C1(
        n258), .Y(n501) );
  OAI222XL U658 ( .A0(n621), .A1(n597), .B0(n724), .B1(n220), .C0(n620), .C1(
        n622), .Y(n577) );
  OAI222XL U659 ( .A0(n130), .A1(n257), .B0(n129), .B1(n1018), .C0(n139), .C1(
        n256), .Y(n969) );
  CLKMX2X2 U660 ( .A(n221), .B(n219), .S0(n246), .Y(n176) );
  OAI221XL U661 ( .A0(n995), .A1(n544), .B0(n543), .B1(n541), .C0(n540), .Y(
        n546) );
  AO21X1 U662 ( .A0(n538), .A1(n537), .B0(n624), .Y(n540) );
  NOR4X1 U663 ( .A(n532), .B(n531), .C(n529), .D(n528), .Y(n543) );
  OAI221XL U664 ( .A0(n995), .A1(n513), .B0(n511), .B1(n541), .C0(n510), .Y(
        n514) );
  AO21X1 U665 ( .A0(n508), .A1(n537), .B0(n620), .Y(n510) );
  NOR4X1 U666 ( .A(n505), .B(n504), .C(n502), .D(n501), .Y(n511) );
  OAI221XL U667 ( .A0(n728), .A1(n269), .B0(n727), .B1(n248), .C0(n726), .Y(
        n736) );
  OA22X1 U668 ( .A0(n232), .A1(n725), .B0(n215), .B1(n724), .Y(n726) );
  MXI2X1 U669 ( .A(n145), .B(n166), .S0(Immediate_SE[8]), .Y(n169) );
  MXI2X1 U670 ( .A(n167), .B(n1018), .S0(n245), .Y(n166) );
  CLKMX2X2 U671 ( .A(n299), .B(n293), .S0(n449), .Y(n450) );
  CLKMX2X2 U672 ( .A(n299), .B(n293), .S0(n385), .Y(n386) );
  CLKMX2X2 U673 ( .A(n299), .B(n293), .S0(n416), .Y(n417) );
  AOI2BB1X1 U674 ( .A0N(n290), .A1N(n944), .B0(n943), .Y(n945) );
  CLKMX2X2 U675 ( .A(n300), .B(n292), .S0(n942), .Y(n944) );
  OR4X1 U676 ( .A(n736), .B(n141), .C(n142), .D(n143), .Y(n742) );
  OAI22XL U677 ( .A0(n256), .A1(n729), .B0(n258), .B1(n329), .Y(n141) );
  OAI22XL U678 ( .A0(n330), .A1(n1018), .B0(n331), .B1(n257), .Y(n142) );
  OR4X1 U679 ( .A(n735), .B(n734), .C(n733), .D(n732), .Y(n143) );
  NAND4X1 U680 ( .A(n477), .B(n475), .C(n474), .D(n472), .Y(n486) );
  OAI222XL U681 ( .A0(n130), .A1(n256), .B0(n158), .B1(n257), .C0(n139), .C1(
        n258), .Y(n378) );
  AOI2BB1X1 U682 ( .A0N(n290), .A1N(n562), .B0(n623), .Y(n563) );
  CLKMX2X2 U683 ( .A(n299), .B(n293), .S0(n561), .Y(n562) );
  AOI2BB1X1 U684 ( .A0N(n290), .A1N(n583), .B0(n582), .Y(n584) );
  CLKMX2X2 U685 ( .A(n299), .B(n293), .S0(n581), .Y(n583) );
  CLKMX2X2 U686 ( .A(n300), .B(n293), .S0(n964), .Y(n966) );
  AOI2BB1X1 U687 ( .A0N(n290), .A1N(n739), .B0(n738), .Y(n740) );
  CLKMX2X2 U688 ( .A(n299), .B(n293), .S0(n737), .Y(n739) );
  CLKMX2X2 U689 ( .A(n299), .B(n293), .S0(n977), .Y(n979) );
  NAND2X1 U690 ( .A(n149), .B(n833), .Y(n830) );
  NAND2X1 U691 ( .A(n149), .B(n808), .Y(n805) );
  NAND2X1 U692 ( .A(n149), .B(n821), .Y(n818) );
  NAND2X1 U693 ( .A(n296), .B(n921), .Y(n918) );
  NAND2X1 U694 ( .A(n149), .B(n237), .Y(n856) );
  NAND2X1 U695 ( .A(n296), .B(n846), .Y(n843) );
  NAND2X1 U696 ( .A(n149), .B(n234), .Y(n906) );
  NAND2X1 U697 ( .A(n149), .B(n236), .Y(n869) );
  NAND2X1 U698 ( .A(n149), .B(n896), .Y(n893) );
  NAND2X1 U699 ( .A(n149), .B(n235), .Y(n881) );
  NAND2X1 U700 ( .A(n149), .B(n943), .Y(n937) );
  NAND2X1 U701 ( .A(n296), .B(n727), .Y(n396) );
  NAND2X1 U702 ( .A(n296), .B(n620), .Y(n496) );
  NAND2X1 U703 ( .A(n296), .B(n624), .Y(n525) );
  NAND2X1 U704 ( .A(n296), .B(n623), .Y(n555) );
  NAND2X1 U705 ( .A(n296), .B(n582), .Y(n572) );
  NAND2X1 U706 ( .A(n296), .B(n606), .Y(n593) );
  NAND2X1 U707 ( .A(n296), .B(n677), .Y(n618) );
  NAND2X1 U708 ( .A(n296), .B(n738), .Y(n722) );
  NAND2X1 U709 ( .A(n149), .B(n257), .Y(n993) );
  MXI4X1 U710 ( .A(n227), .B(n219), .C(n221), .D(n1018), .S0(n245), .S1(n246), 
        .Y(n144) );
  MXI4X1 U711 ( .A(n201), .B(n222), .C(n223), .D(n1018), .S0(n245), .S1(n246), 
        .Y(n146) );
  CLKMX2X2 U712 ( .A(n535), .B(n294), .S0(n534), .Y(n538) );
  CLKMX2X2 U713 ( .A(n535), .B(n291), .S0(n507), .Y(n508) );
  OR4X1 U714 ( .A(n580), .B(n579), .C(n578), .D(n577), .Y(n586) );
  OAI222XL U715 ( .A0(n139), .A1(n623), .B0(n624), .B1(n130), .C0(n582), .C1(
        n177), .Y(n578) );
  OAI222XL U716 ( .A0(n727), .A1(n575), .B0(n728), .B1(n574), .C0(n725), .C1(
        n596), .Y(n580) );
  OAI221XL U717 ( .A0(n268), .A1(n1018), .B0(n257), .B1(n269), .C0(n576), .Y(
        n579) );
  CLKMX2X2 U718 ( .A(n210), .B(n209), .S0(n246), .Y(n172) );
  CLKMX2X2 U719 ( .A(n223), .B(n222), .S0(n246), .Y(n167) );
  CLKMX2X2 U720 ( .A(n299), .B(n293), .S0(n767), .Y(n769) );
  CLKMX2X2 U721 ( .A(n299), .B(n292), .S0(n794), .Y(n796) );
  CLKMX2X2 U722 ( .A(n300), .B(n292), .S0(n820), .Y(n822) );
  CLKMX2X2 U723 ( .A(n300), .B(n292), .S0(n895), .Y(n897) );
  AOI2BB1X1 U724 ( .A0N(n290), .A1N(n678), .B0(n677), .Y(n712) );
  CLKMX2X2 U725 ( .A(n299), .B(n293), .S0(n676), .Y(n678) );
  CLKMX2X2 U726 ( .A(n299), .B(n293), .S0(n754), .Y(n756) );
  CLKMX2X2 U727 ( .A(n300), .B(n292), .S0(n858), .Y(n859) );
  AOI2BB1X1 U728 ( .A0N(n1000), .A1N(n401), .B0(n727), .Y(n402) );
  CLKMX2X2 U729 ( .A(n299), .B(n293), .S0(n400), .Y(n401) );
  AOI2BB1X1 U730 ( .A0N(n290), .A1N(n607), .B0(n606), .Y(n608) );
  CLKMX2X2 U731 ( .A(n299), .B(n293), .S0(n605), .Y(n607) );
  AOI2BB1X1 U732 ( .A0N(n1000), .A1N(n999), .B0(n257), .Y(n1001) );
  CLKMX2X2 U733 ( .A(n299), .B(n293), .S0(n996), .Y(n999) );
  CLKMX2X2 U734 ( .A(n300), .B(n292), .S0(n883), .Y(n884) );
  CLKMX2X2 U735 ( .A(n300), .B(n293), .S0(n953), .Y(n955) );
  CLKMX2X2 U736 ( .A(n300), .B(n292), .S0(n845), .Y(n847) );
  CLKMX2X2 U737 ( .A(n300), .B(n292), .S0(n871), .Y(n872) );
  CLKMX2X2 U738 ( .A(n300), .B(n292), .S0(n920), .Y(n922) );
  CLKMX2X2 U739 ( .A(n299), .B(n293), .S0(n780), .Y(n782) );
  CLKMX2X2 U740 ( .A(n300), .B(n292), .S0(n807), .Y(n809) );
  CLKMX2X2 U741 ( .A(n300), .B(n292), .S0(n832), .Y(n834) );
  CLKMX2X2 U742 ( .A(n300), .B(n292), .S0(n908), .Y(n909) );
  AND2X2 U743 ( .A(n1012), .B(n326), .Y(n148) );
  AND2X2 U744 ( .A(n161), .B(n327), .Y(n149) );
  AND2X2 U745 ( .A(n159), .B(n325), .Y(n150) );
  AND2X2 U746 ( .A(n160), .B(n332), .Y(n151) );
  AND2X2 U747 ( .A(n1008), .B(n332), .Y(n152) );
  NAND2X1 U748 ( .A(n153), .B(n940), .Y(n383) );
  AOI21X1 U749 ( .A0(n350), .A1(n348), .B0(n317), .Y(n330) );
  CLKINVX1 U750 ( .A(n382), .Y(n1020) );
  NAND2X1 U751 ( .A(n349), .B(n354), .Y(n248) );
  AND2X2 U752 ( .A(n384), .B(n333), .Y(n1000) );
  OAI21XL U753 ( .A0(n383), .A1(n177), .B0(n382), .Y(n384) );
  NAND2X1 U754 ( .A(n350), .B(n354), .Y(n269) );
  NAND2X1 U755 ( .A(n349), .B(n351), .Y(n329) );
  CLKINVX1 U756 ( .A(n1009), .Y(n1016) );
  NAND2X1 U757 ( .A(n348), .B(n349), .Y(n331) );
  AND2X2 U758 ( .A(n155), .B(n1014), .Y(n153) );
  AND2X2 U759 ( .A(n350), .B(n351), .Y(n313) );
  CLKBUFX3 U760 ( .A(n337), .Y(n334) );
  CLKBUFX3 U761 ( .A(n337), .Y(n335) );
  CLKBUFX3 U762 ( .A(n337), .Y(n336) );
  NAND2X2 U763 ( .A(n358), .B(n353), .Y(n139) );
  NAND2X2 U764 ( .A(n359), .B(n354), .Y(n130) );
  NAND2X1 U765 ( .A(n351), .B(n358), .Y(n220) );
  CLKBUFX3 U766 ( .A(n451), .Y(n306) );
  CLKBUFX3 U767 ( .A(n451), .Y(n305) );
  CLKBUFX3 U768 ( .A(n453), .Y(n303) );
  CLKBUFX3 U769 ( .A(n455), .Y(n302) );
  CLKBUFX3 U770 ( .A(n455), .Y(n301) );
  CLKBUFX3 U771 ( .A(n453), .Y(n304) );
  CLKBUFX3 U772 ( .A(n339), .Y(n340) );
  CLKMX2X2 U773 ( .A(n938), .B(n937), .S0(n942), .Y(n949) );
  AOI211X1 U774 ( .A0(N493), .A1(n284), .B0(n946), .C0(n945), .Y(n947) );
  MXI2XL U775 ( .A(n108), .B(ALUData2[15]), .S0(n249), .Y(n226) );
  MXI2XL U776 ( .A(ALUData2[12]), .B(ALUData2[13]), .S0(n249), .Y(n193) );
  MXI2XL U777 ( .A(n134), .B(ALUData2[12]), .S0(n249), .Y(n196) );
  MXI2XL U778 ( .A(ALUData2[10]), .B(n134), .S0(n249), .Y(n201) );
  MXI2XL U779 ( .A(ALUData2[13]), .B(n108), .S0(n249), .Y(n190) );
  NAND2X1 U780 ( .A(n320), .B(ALUresult[30]), .Y(n1006) );
  NAND2X1 U781 ( .A(n320), .B(ALUresult[27]), .Y(n392) );
  NAND2X1 U782 ( .A(n320), .B(ALUresult[29]), .Y(n988) );
  CLKMX2X2 U783 ( .A(n976), .B(n975), .S0(n977), .Y(n987) );
  NOR4X1 U784 ( .A(n985), .B(n984), .C(n109), .D(n983), .Y(n986) );
  NAND2X1 U785 ( .A(n321), .B(ALUresult[19]), .Y(n589) );
  AOI211X1 U786 ( .A0(n284), .A1(n586), .B0(n585), .C0(n584), .Y(n587) );
  NAND2X1 U787 ( .A(n321), .B(n430), .Y(n463) );
  NOR4X1 U788 ( .A(n459), .B(n457), .C(n456), .D(n452), .Y(n460) );
  NAND2X1 U789 ( .A(n321), .B(n411), .Y(n424) );
  NOR4X1 U790 ( .A(n421), .B(n420), .C(n419), .D(n418), .Y(n422) );
  NAND2X1 U791 ( .A(n321), .B(ALUresult[23]), .Y(n490) );
  AOI211X1 U792 ( .A0(n284), .A1(n486), .B0(n484), .C0(n483), .Y(n487) );
  NAND2X1 U793 ( .A(n320), .B(ALUresult[15]), .Y(n960) );
  CLKMX2X2 U794 ( .A(n952), .B(n951), .S0(n953), .Y(n959) );
  NAND2X1 U795 ( .A(n321), .B(ALUresult[14]), .Y(n761) );
  CLKMX2X2 U796 ( .A(n753), .B(n752), .S0(n754), .Y(n760) );
  NAND2X1 U797 ( .A(n321), .B(ALUresult[13]), .Y(n774) );
  CLKMX2X2 U798 ( .A(n766), .B(n765), .S0(n767), .Y(n773) );
  NAND2X1 U799 ( .A(n321), .B(ALUresult[12]), .Y(n787) );
  CLKMX2X2 U800 ( .A(n779), .B(n778), .S0(n780), .Y(n786) );
  NAND2X1 U801 ( .A(n320), .B(ALUresult[11]), .Y(n801) );
  CLKMX2X2 U802 ( .A(n793), .B(n792), .S0(n794), .Y(n800) );
  NAND2X1 U803 ( .A(n321), .B(ALUresult[10]), .Y(n814) );
  CLKMX2X2 U804 ( .A(n806), .B(n805), .S0(n807), .Y(n813) );
  NAND2X1 U805 ( .A(n321), .B(ALUresult[9]), .Y(n827) );
  CLKMX2X2 U806 ( .A(n819), .B(n818), .S0(n820), .Y(n826) );
  NAND2X1 U807 ( .A(n320), .B(ALUresult[8]), .Y(n839) );
  CLKMX2X2 U808 ( .A(n831), .B(n830), .S0(n832), .Y(n838) );
  NAND2X1 U809 ( .A(n321), .B(ALUresult[7]), .Y(n852) );
  CLKMX2X2 U810 ( .A(n844), .B(n843), .S0(n845), .Y(n851) );
  NAND2X1 U811 ( .A(n320), .B(ALUresult[6]), .Y(n864) );
  CLKMX2X2 U812 ( .A(n857), .B(n856), .S0(n858), .Y(n863) );
  NAND2X1 U813 ( .A(n320), .B(ALUresult[5]), .Y(n877) );
  CLKMX2X2 U814 ( .A(n870), .B(n869), .S0(n871), .Y(n876) );
  NAND2X1 U815 ( .A(n320), .B(ALUresult[4]), .Y(n889) );
  CLKMX2X2 U816 ( .A(n882), .B(n881), .S0(n883), .Y(n888) );
  NAND2X1 U817 ( .A(n320), .B(ALUresult[3]), .Y(n902) );
  CLKMX2X2 U818 ( .A(n894), .B(n893), .S0(n895), .Y(n901) );
  NAND2X1 U819 ( .A(n320), .B(ALUresult[2]), .Y(n914) );
  CLKMX2X2 U820 ( .A(n907), .B(n906), .S0(n908), .Y(n913) );
  NAND4BX1 U821 ( .AN(n928), .B(n927), .C(n926), .D(n925), .Y(
        next_ALUresult[1]) );
  NAND2X1 U822 ( .A(n320), .B(ALUresult[1]), .Y(n927) );
  CLKMX2X2 U823 ( .A(n919), .B(n918), .S0(n920), .Y(n926) );
  AO22X1 U824 ( .A0(N333), .A1(n151), .B0(N205), .B1(n152), .Y(n928) );
  NAND2X1 U825 ( .A(n321), .B(ALUresult[17]), .Y(n717) );
  CLKMX2X2 U826 ( .A(n619), .B(n618), .S0(n676), .Y(n716) );
  AOI211X1 U827 ( .A0(n284), .A1(n714), .B0(n713), .C0(n712), .Y(n715) );
  NAND2X1 U828 ( .A(n321), .B(ALUresult[18]), .Y(n613) );
  CLKMX2X2 U829 ( .A(n594), .B(n593), .S0(n605), .Y(n612) );
  AOI211X1 U830 ( .A0(n284), .A1(n610), .B0(n609), .C0(n608), .Y(n611) );
  NAND2X1 U831 ( .A(n321), .B(ALUresult[20]), .Y(n568) );
  AOI211X1 U832 ( .A0(n284), .A1(n565), .B0(n564), .C0(n563), .Y(n566) );
  NAND2X1 U833 ( .A(n321), .B(ALUresult[16]), .Y(n745) );
  CLKMX2X2 U834 ( .A(n723), .B(n722), .S0(n737), .Y(n744) );
  AOI211X1 U835 ( .A0(n284), .A1(n742), .B0(n741), .C0(n740), .Y(n743) );
  NAND2X1 U836 ( .A(n321), .B(ALUresult[26]), .Y(n407) );
  AOI211X1 U837 ( .A0(n284), .A1(n404), .B0(n403), .C0(n402), .Y(n405) );
  NAND2X1 U838 ( .A(n321), .B(ALUresult[21]), .Y(n550) );
  NAND2X1 U839 ( .A(n321), .B(ALUresult[22]), .Y(n519) );
  NAND2X1 U840 ( .A(n320), .B(ALUresult[28]), .Y(n972) );
  AOI211X1 U841 ( .A0(n284), .A1(n969), .B0(n968), .C0(n967), .Y(n970) );
  CLKINVX1 U842 ( .A(WBData[11]), .Y(n1063) );
  MXI2X1 U843 ( .A(n206), .B(n202), .S0(Immediate_SE[7]), .Y(N493) );
  MX3XL U844 ( .A(n233), .B(n176), .C(n230), .S0(Immediate_SE[10]), .S1(
        Immediate_SE[8]), .Y(n206) );
  MXI3XL U845 ( .A(n5), .B(ALUData2[1]), .C(n238), .S0(Immediate_SE[6]), .S1(
        Immediate_SE[9]), .Y(n233) );
  CLKINVX1 U846 ( .A(n227), .Y(n238) );
  MXI3X1 U847 ( .A(n203), .B(n241), .C(n125), .S0(Immediate_SE[10]), .S1(
        Immediate_SE[8]), .Y(n205) );
  MXI3X1 U848 ( .A(n236), .B(n237), .C(n190), .S0(n249), .S1(n246), .Y(n189)
         );
  INVXL U849 ( .A(ALUData2[6]), .Y(n237) );
  MXI2XL U850 ( .A(ALUData2[7]), .B(ALUData2[8]), .S0(n249), .Y(n228) );
  MXI2XL U851 ( .A(ALUData2[6]), .B(ALUData2[7]), .S0(n249), .Y(n229) );
  INVXL U852 ( .A(ALUData2[12]), .Y(n781) );
  INVXL U853 ( .A(ALUData2[8]), .Y(n833) );
  INVXL U854 ( .A(ALUData2[10]), .Y(n808) );
  INVXL U855 ( .A(ALUData2[13]), .Y(n768) );
  INVXL U856 ( .A(n134), .Y(n795) );
  INVXL U857 ( .A(ALUData2[9]), .Y(n821) );
  INVXL U858 ( .A(ALUData2[1]), .Y(n921) );
  INVXL U859 ( .A(ALUData2[15]), .Y(n954) );
  INVXL U860 ( .A(ALUData2[14]), .Y(n755) );
  INVXL U861 ( .A(ALUData2[7]), .Y(n846) );
  INVXL U862 ( .A(n5), .Y(n943) );
  INVXL U863 ( .A(ALUData1[13]), .Y(n767) );
  INVXL U864 ( .A(ALUData1[11]), .Y(n794) );
  INVXL U865 ( .A(n702), .Y(n820) );
  INVXL U866 ( .A(ALUData1[3]), .Y(n895) );
  INVXL U867 ( .A(ALUData1[17]), .Y(n676) );
  INVXL U868 ( .A(ALUData1[24]), .Y(n449) );
  INVXL U869 ( .A(ALUData1[20]), .Y(n561) );
  INVXL U870 ( .A(ALUData1[14]), .Y(n754) );
  INVXL U871 ( .A(ALUData1[6]), .Y(n858) );
  INVXL U872 ( .A(ALUData1[18]), .Y(n605) );
  INVXL U873 ( .A(ALUData1[4]), .Y(n883) );
  INVXL U874 ( .A(ALUData1[19]), .Y(n581) );
  INVXL U875 ( .A(ALUData1[21]), .Y(n534) );
  INVXL U876 ( .A(ALUData1[25]), .Y(n416) );
  INVXL U877 ( .A(ALUData1[15]), .Y(n953) );
  INVXL U878 ( .A(ALUData1[7]), .Y(n845) );
  INVXL U879 ( .A(ALUData1[5]), .Y(n871) );
  INVXL U880 ( .A(ALUData1[1]), .Y(n920) );
  INVXL U881 ( .A(ALUData1[12]), .Y(n780) );
  INVXL U882 ( .A(ALUData1[10]), .Y(n807) );
  INVXL U883 ( .A(ALUData1[8]), .Y(n832) );
  INVXL U884 ( .A(ALUData1[2]), .Y(n908) );
  MXI2XL U885 ( .A(ALUData2[9]), .B(ALUData2[10]), .S0(n249), .Y(n204) );
  OAI221XL U886 ( .A0(n130), .A1(n258), .B0(n139), .B1(n728), .C0(n399), .Y(
        n404) );
  AOI222XL U887 ( .A0(n253), .A1(n1111), .B0(n251), .B1(n398), .C0(n252), .C1(
        n731), .Y(n399) );
  AOI222XL U888 ( .A0(n1115), .A1(n259), .B0(n625), .B1(n254), .C0(n1112), 
        .C1(n255), .Y(n559) );
  NOR4X1 U889 ( .A(n630), .B(n629), .C(n628), .D(n627), .Y(n631) );
  AO22X1 U890 ( .A0(n1112), .A1(n261), .B0(n260), .B1(n625), .Y(n630) );
  AO22X1 U891 ( .A0(n259), .A1(n626), .B0(n255), .B1(n1109), .Y(n629) );
  AO22X1 U892 ( .A0(n1108), .A1(n254), .B0(n253), .B1(n1110), .Y(n628) );
  AOI31X1 U893 ( .A0(n440), .A1(n438), .A2(n437), .B0(n541), .Y(n457) );
  OA22X1 U894 ( .A0(n186), .A1(n257), .B0(n256), .B1(n220), .Y(n440) );
  AOI222XL U895 ( .A0(n1114), .A1(n261), .B0(n1113), .B1(n259), .C0(n260), 
        .C1(n981), .Y(n437) );
  OA22X1 U896 ( .A0(n258), .A1(n597), .B0(n728), .B1(n622), .Y(n438) );
  CLKINVX1 U897 ( .A(WBData[19]), .Y(n1055) );
  CLKINVX1 U898 ( .A(WBData[14]), .Y(n1060) );
  CLKINVX1 U899 ( .A(WBData[23]), .Y(n1051) );
  CLKINVX1 U900 ( .A(WBData[16]), .Y(n1058) );
  CLKINVX1 U901 ( .A(WBData[17]), .Y(n1057) );
  CLKINVX1 U902 ( .A(WBData[26]), .Y(n1048) );
  CLKINVX1 U903 ( .A(WBData[24]), .Y(n1050) );
  CLKINVX1 U904 ( .A(WBData[27]), .Y(n1047) );
  CLKINVX1 U905 ( .A(WBData[13]), .Y(n1061) );
  CLKINVX1 U906 ( .A(WBData[18]), .Y(n1056) );
  CLKINVX1 U907 ( .A(WBData[30]), .Y(n1044) );
  CLKINVX1 U908 ( .A(WBData[31]), .Y(n1043) );
  CLKINVX1 U909 ( .A(WBData[21]), .Y(n1053) );
  CLKINVX1 U910 ( .A(WBData[22]), .Y(n1052) );
  CLKINVX1 U911 ( .A(WBData[20]), .Y(n1054) );
  CLKINVX1 U912 ( .A(WBData[1]), .Y(n1039) );
  CLKINVX1 U913 ( .A(WBData[0]), .Y(n1035) );
  CLKINVX1 U914 ( .A(WBData[4]), .Y(n1070) );
  CLKINVX1 U915 ( .A(WBData[9]), .Y(n1065) );
  AOI2BB1X1 U916 ( .A0N(n415), .A1N(n414), .B0(n541), .Y(n420) );
  OAI222XL U917 ( .A0(n256), .A1(n597), .B0(n257), .B1(n220), .C0(n158), .C1(
        n258), .Y(n414) );
  NAND4X1 U918 ( .A(n604), .B(n603), .C(n602), .D(n601), .Y(n610) );
  AOI222XL U919 ( .A0(n260), .A1(n1112), .B0(n255), .B1(n626), .C0(n259), .C1(
        n625), .Y(n602) );
  OA22X1 U920 ( .A0(n256), .A1(n269), .B0(n258), .B1(n248), .Y(n603) );
  OA22X1 U921 ( .A0(n1018), .A1(n595), .B0(n257), .B1(n329), .Y(n604) );
  NAND4X1 U922 ( .A(n675), .B(n674), .C(n636), .D(n631), .Y(n714) );
  AOI222XL U923 ( .A0(n1114), .A1(n270), .B0(n1113), .B1(n266), .C0(n267), 
        .C1(n981), .Y(n636) );
  OA22X1 U924 ( .A0(n157), .A1(n624), .B0(n623), .B1(n622), .Y(n674) );
  OA22X1 U925 ( .A0(n186), .A1(n621), .B0(n620), .B1(n220), .Y(n675) );
  NAND4X1 U926 ( .A(n560), .B(n559), .C(n558), .D(n557), .Y(n565) );
  AOI222XL U927 ( .A0(n626), .A1(n253), .B0(n247), .B1(n251), .C0(n1109), .C1(
        n252), .Y(n560) );
  AOI222XL U928 ( .A0(n1114), .A1(n265), .B0(n1113), .B1(n263), .C0(n264), 
        .C1(n981), .Y(n557) );
  AOI222XL U929 ( .A0(n1111), .A1(n262), .B0(n730), .B1(n260), .C0(n731), .C1(
        n261), .Y(n558) );
  AOI2BB1XL U930 ( .A0N(ALUData2[12]), .A1N(n291), .B0(n288), .Y(n779) );
  AOI2BB1XL U931 ( .A0N(ALUData2[8]), .A1N(n992), .B0(n289), .Y(n831) );
  AOI2BB1XL U932 ( .A0N(ALUData2[10]), .A1N(n294), .B0(n288), .Y(n806) );
  AOI2BB1XL U933 ( .A0N(ALUData2[13]), .A1N(n291), .B0(n288), .Y(n766) );
  AOI2BB1XL U934 ( .A0N(n134), .A1N(n291), .B0(n288), .Y(n793) );
  AOI2BB1XL U935 ( .A0N(ALUData2[9]), .A1N(n291), .B0(n288), .Y(n819) );
  AOI2BB1XL U936 ( .A0N(ALUData2[1]), .A1N(n992), .B0(n288), .Y(n919) );
  AOI2BB1XL U937 ( .A0N(ALUData2[6]), .A1N(n294), .B0(n290), .Y(n857) );
  AOI2BB1XL U938 ( .A0N(ALUData2[15]), .A1N(n291), .B0(n288), .Y(n952) );
  AOI2BB1XL U939 ( .A0N(n108), .A1N(n291), .B0(n288), .Y(n753) );
  AOI2BB1XL U940 ( .A0N(ALUData2[7]), .A1N(n992), .B0(n290), .Y(n844) );
  AOI2BB1XL U941 ( .A0N(ALUData2[2]), .A1N(n291), .B0(n288), .Y(n907) );
  AOI2BB1XL U942 ( .A0N(ALUData2[5]), .A1N(n291), .B0(n288), .Y(n870) );
  AOI2BB1XL U943 ( .A0N(ALUData2[3]), .A1N(n992), .B0(n288), .Y(n894) );
  AOI2BB1XL U944 ( .A0N(ALUData2[4]), .A1N(n992), .B0(n288), .Y(n882) );
  AOI2BB1XL U945 ( .A0N(n5), .A1N(n291), .B0(n290), .Y(n938) );
  CLKINVX1 U946 ( .A(n164), .Y(n243) );
  AO22X1 U947 ( .A0(n481), .A1(n262), .B0(n197), .B1(n980), .Y(n483) );
  NAND2X1 U948 ( .A(n480), .B(n537), .Y(n481) );
  CLKMX2X2 U949 ( .A(n535), .B(n294), .S0(n478), .Y(n480) );
  AO22X1 U950 ( .A0(n265), .A1(n731), .B0(n264), .B1(n730), .Y(n733) );
  CLKBUFX3 U951 ( .A(n965), .Y(n258) );
  CLKINVX1 U952 ( .A(n254), .Y(n965) );
  CLKBUFX3 U953 ( .A(n978), .Y(n256) );
  CLKINVX1 U954 ( .A(n253), .Y(n978) );
  AND3X2 U955 ( .A(n600), .B(n599), .C(n598), .Y(n601) );
  AOI222XL U956 ( .A0(n1114), .A1(n267), .B0(n1113), .B1(n265), .C0(n266), 
        .C1(n981), .Y(n598) );
  OA22X1 U957 ( .A0(n620), .A1(n597), .B0(n624), .B1(n622), .Y(n599) );
  OA22X1 U958 ( .A0(n724), .A1(n596), .B0(n621), .B1(n220), .Y(n600) );
  AO22X1 U959 ( .A0(n1113), .A1(n267), .B0(n1111), .B1(n266), .Y(n734) );
  CLKMX2X2 U960 ( .A(n1017), .B(n1016), .S0(n1015), .Y(n1019) );
  AND2X2 U961 ( .A(n1014), .B(n1013), .Y(n1017) );
  AO22X1 U962 ( .A0(n264), .A1(n1114), .B0(n263), .B1(n981), .Y(n532) );
  AO22X1 U963 ( .A0(n263), .A1(n1114), .B0(n262), .B1(n981), .Y(n505) );
  NAND3BX1 U964 ( .AN(n322), .B(n1014), .C(n1013), .Y(n535) );
  CLKINVX1 U965 ( .A(n939), .Y(n1014) );
  CLKINVX1 U966 ( .A(n373), .Y(n1008) );
  NAND2X1 U967 ( .A(n439), .B(n1119), .Y(n434) );
  CLKINVX1 U968 ( .A(stall), .Y(n337) );
  CLKINVX1 U969 ( .A(n379), .Y(n1012) );
  CLKBUFX3 U970 ( .A(rst), .Y(n339) );
  CLKBUFX3 U971 ( .A(rst), .Y(n338) );
  CLKMX2X2 U972 ( .A(n941), .B(n1148), .S0(n320), .Y(n948) );
  NAND4X1 U973 ( .A(N524), .B(n155), .C(n940), .D(n939), .Y(n941) );
  CLKINVX1 U974 ( .A(Immediate_SE[5]), .Y(n867) );
  OA22X1 U975 ( .A0(n1070), .A1(n282), .B0(n1105), .B1(n279), .Y(n879) );
  OA22X1 U976 ( .A0(n282), .A1(n1035), .B0(n278), .B1(n1036), .Y(n934) );
  NAND2X1 U977 ( .A(RData1[11]), .B(n6), .Y(n788) );
  NAND2X1 U978 ( .A(RData1[9]), .B(n6), .Y(n815) );
  NAND2X1 U979 ( .A(RData1[20]), .B(n6), .Y(n552) );
  NAND2X1 U980 ( .A(RData1[6]), .B(n6), .Y(n853) );
  NAND2X1 U981 ( .A(RData1[22]), .B(n6), .Y(n493) );
  NAND2X1 U982 ( .A(RData1[7]), .B(n6), .Y(n840) );
  OAI221XL U983 ( .A0(n1043), .A1(n281), .B0(n1078), .B1(n280), .C0(n360), .Y(
        ALUData2[31]) );
  AOI2BB2X1 U984 ( .B0(Immediate_SE[31]), .B1(n789), .A0N(n679), .A1N(n283), 
        .Y(n360) );
  NAND2X1 U985 ( .A(RData1[25]), .B(n6), .Y(n409) );
  OAI221XL U986 ( .A0(n1048), .A1(n282), .B0(n1083), .B1(n280), .C0(n395), .Y(
        ALUData2[26]) );
  AOI2BB2X1 U987 ( .B0(Immediate_SE[26]), .B1(n789), .A0N(n684), .A1N(n283), 
        .Y(n395) );
  OAI221XL U988 ( .A0(n1047), .A1(n282), .B0(n1082), .B1(n278), .C0(n371), .Y(
        ALUData2[27]) );
  AOI2BB2X1 U989 ( .B0(Immediate_SE[27]), .B1(n789), .A0N(n683), .A1N(n283), 
        .Y(n371) );
  BUFX4 U990 ( .A(ALUData2[25]), .Y(n260) );
  OAI221XL U991 ( .A0(n1049), .A1(n282), .B0(n1084), .B1(n280), .C0(n410), .Y(
        ALUData2[25]) );
  AOI2BB2X1 U992 ( .B0(Immediate_SE[25]), .B1(n789), .A0N(n685), .A1N(n283), 
        .Y(n410) );
  OAI221XL U993 ( .A0(n1044), .A1(n282), .B0(n1079), .B1(n278), .C0(n364), .Y(
        ALUData2[30]) );
  AOI2BB2X1 U994 ( .B0(Immediate_SE[30]), .B1(n789), .A0N(n680), .A1N(n283), 
        .Y(n364) );
  BUFX4 U995 ( .A(ALUData2[24]), .Y(n261) );
  OAI221XL U996 ( .A0(n1050), .A1(n282), .B0(n1085), .B1(n280), .C0(n427), .Y(
        ALUData2[24]) );
  AOI2BB2X1 U997 ( .B0(Immediate_SE[24]), .B1(n789), .A0N(n686), .A1N(n283), 
        .Y(n427) );
  OAI221XL U998 ( .A0(n1045), .A1(n282), .B0(n1080), .B1(n278), .C0(n367), .Y(
        ALUData2[29]) );
  AOI2BB2X1 U999 ( .B0(Immediate_SE[29]), .B1(n789), .A0N(n681), .A1N(n283), 
        .Y(n367) );
  OAI221XL U1000 ( .A0(n1051), .A1(n282), .B0(n1086), .B1(n278), .C0(n468), 
        .Y(ALUData2[23]) );
  AOI2BB2X1 U1001 ( .B0(Immediate_SE[23]), .B1(n789), .A0N(n687), .A1N(n283), 
        .Y(n468) );
  OAI221XL U1002 ( .A0(n1052), .A1(n281), .B0(n1087), .B1(n278), .C0(n495), 
        .Y(ALUData2[22]) );
  AOI2BB2X1 U1003 ( .B0(Immediate_SE[22]), .B1(n789), .A0N(n688), .A1N(n283), 
        .Y(n495) );
  OAI221XL U1004 ( .A0(n1046), .A1(n282), .B0(n1081), .B1(n278), .C0(n368), 
        .Y(ALUData2[28]) );
  AOI2BB2X1 U1005 ( .B0(Immediate_SE[28]), .B1(n789), .A0N(n682), .A1N(n283), 
        .Y(n368) );
  BUFX4 U1006 ( .A(ALUData2[20]), .Y(n265) );
  OAI221XL U1007 ( .A0(n1054), .A1(n281), .B0(n1089), .B1(n280), .C0(n553), 
        .Y(ALUData2[20]) );
  AOI2BB2X1 U1008 ( .B0(Immediate_SE[20]), .B1(n789), .A0N(n690), .A1N(n283), 
        .Y(n553) );
  OAI221XL U1009 ( .A0(n1056), .A1(n281), .B0(n1091), .B1(n280), .C0(n592), 
        .Y(ALUData2[18]) );
  AOI2BB2X1 U1010 ( .B0(Immediate_SE[18]), .B1(n789), .A0N(n692), .A1N(n283), 
        .Y(n592) );
  OAI221XL U1011 ( .A0(n1055), .A1(n281), .B0(n1090), .B1(n280), .C0(n571), 
        .Y(ALUData2[19]) );
  AOI2BB2X1 U1012 ( .B0(Immediate_SE[19]), .B1(n789), .A0N(n691), .A1N(n283), 
        .Y(n571) );
  OAI221XL U1013 ( .A0(n1053), .A1(n281), .B0(n1088), .B1(n280), .C0(n523), 
        .Y(ALUData2[21]) );
  AOI2BB2X1 U1014 ( .B0(Immediate_SE[21]), .B1(n789), .A0N(n689), .A1N(n283), 
        .Y(n523) );
  BUFX4 U1015 ( .A(ALUData2[17]), .Y(n270) );
  OAI221XL U1016 ( .A0(n1057), .A1(n281), .B0(n1092), .B1(n280), .C0(n616), 
        .Y(ALUData2[17]) );
  AOI2BB2X1 U1017 ( .B0(Immediate_SE[17]), .B1(n789), .A0N(n693), .A1N(n283), 
        .Y(n616) );
  CLKBUFX3 U1018 ( .A(ALUData2[16]), .Y(n271) );
  OAI221XL U1019 ( .A0(n1058), .A1(n281), .B0(n1093), .B1(n280), .C0(n720), 
        .Y(ALUData2[16]) );
  AOI2BB2X1 U1020 ( .B0(Immediate_SE[16]), .B1(n789), .A0N(n694), .A1N(n283), 
        .Y(n720) );
  CLKINVX1 U1021 ( .A(RData2[11]), .Y(n1098) );
  CLKINVX1 U1022 ( .A(ID_EX[2]), .Y(n372) );
  NAND2X1 U1023 ( .A(n441), .B(ID_EX[2]), .Y(n381) );
  NAND4X1 U1024 ( .A(n1117), .B(n1116), .C(n1120), .D(n442), .Y(n441) );
  NAND2X1 U1025 ( .A(n446), .B(n447), .Y(n939) );
  XOR2X1 U1026 ( .A(ID_EX[2]), .B(ID_EX[1]), .Y(n446) );
  OAI21XL U1027 ( .A0(n448), .A1(n372), .B0(n1042), .Y(n447) );
  CLKINVX1 U1028 ( .A(ID_EX[3]), .Y(n1042) );
  NAND4BX1 U1029 ( .AN(ID_EX[1]), .B(ID_EX[2]), .C(n429), .D(n1042), .Y(n428)
         );
  AOI2BB2X1 U1030 ( .B0(n434), .B1(n435), .A0N(n1118), .A1N(n1117), .Y(n433)
         );
  CLKINVX1 U1031 ( .A(RData2[28]), .Y(n1081) );
  CLKINVX1 U1032 ( .A(RData2[19]), .Y(n1090) );
  CLKINVX1 U1033 ( .A(RData2[17]), .Y(n1092) );
  CLKINVX1 U1034 ( .A(RData2[18]), .Y(n1091) );
  CLKINVX1 U1035 ( .A(RData2[27]), .Y(n1082) );
  CLKINVX1 U1036 ( .A(RData2[26]), .Y(n1083) );
  CLKINVX1 U1037 ( .A(RData2[23]), .Y(n1086) );
  CLKINVX1 U1038 ( .A(RData2[25]), .Y(n1084) );
  CLKINVX1 U1039 ( .A(RData2[24]), .Y(n1085) );
  CLKINVX1 U1040 ( .A(RData2[22]), .Y(n1087) );
  CLKINVX1 U1041 ( .A(RData2[21]), .Y(n1088) );
  CLKINVX1 U1042 ( .A(RData2[20]), .Y(n1089) );
  CLKINVX1 U1043 ( .A(RData2[31]), .Y(n1078) );
  CLKINVX1 U1044 ( .A(RData2[29]), .Y(n1080) );
  CLKINVX1 U1045 ( .A(RData2[30]), .Y(n1079) );
  OA21XL U1046 ( .A0(n1118), .A1(Immediate_SE[1]), .B0(Immediate_SE[5]), .Y(
        n448) );
  OAI221XL U1047 ( .A0(n305), .A1(n1040), .B0(n304), .B1(n1039), .C0(n1038), 
        .Y(n660) );
  OAI221XL U1048 ( .A0(n306), .A1(n1036), .B0(n304), .B1(n1035), .C0(n1034), 
        .Y(n668) );
  OA22X1 U1049 ( .A0(n301), .A1(n1149), .B0(n333), .B1(n905), .Y(n1034) );
  OAI221XL U1050 ( .A0(n1090), .A1(n306), .B0(n1055), .B1(n304), .C0(n454), 
        .Y(n637) );
  AOI2BB2XL U1051 ( .B0(n320), .B1(MEMWriteData[19]), .A0N(n302), .A1N(n691), 
        .Y(n454) );
  OAI221XL U1052 ( .A0(n1088), .A1(n305), .B0(n1053), .B1(n304), .C0(n458), 
        .Y(n638) );
  AOI2BB2XL U1053 ( .B0(n319), .B1(MEMWriteData[21]), .A0N(n302), .A1N(n689), 
        .Y(n458) );
  OAI221XL U1054 ( .A0(n1087), .A1(n451), .B0(n1052), .B1(n304), .C0(n461), 
        .Y(n639) );
  AOI2BB2XL U1055 ( .B0(n319), .B1(MEMWriteData[22]), .A0N(n302), .A1N(n688), 
        .Y(n461) );
  OAI221XL U1056 ( .A0(n1086), .A1(n451), .B0(n1051), .B1(n304), .C0(n464), 
        .Y(n640) );
  AOI2BB2XL U1057 ( .B0(n319), .B1(MEMWriteData[23]), .A0N(n302), .A1N(n687), 
        .Y(n464) );
  OAI221XL U1058 ( .A0(n1085), .A1(n306), .B0(n1050), .B1(n304), .C0(n467), 
        .Y(n641) );
  AOI2BB2XL U1059 ( .B0(n319), .B1(MEMWriteData[24]), .A0N(n302), .A1N(n686), 
        .Y(n467) );
  OAI221XL U1060 ( .A0(n1084), .A1(n306), .B0(n1049), .B1(n304), .C0(n470), 
        .Y(n642) );
  AOI2BB2XL U1061 ( .B0(n319), .B1(MEMWriteData[25]), .A0N(n302), .A1N(n685), 
        .Y(n470) );
  OAI221XL U1062 ( .A0(n1083), .A1(n306), .B0(n1048), .B1(n303), .C0(n473), 
        .Y(n643) );
  AOI2BB2XL U1063 ( .B0(n319), .B1(MEMWriteData[26]), .A0N(n302), .A1N(n684), 
        .Y(n473) );
  OAI221XL U1064 ( .A0(n1082), .A1(n306), .B0(n1047), .B1(n303), .C0(n476), 
        .Y(n644) );
  OA22X1 U1065 ( .A0(n333), .A1(n1143), .B0(n301), .B1(n683), .Y(n476) );
  OAI221XL U1066 ( .A0(n1081), .A1(n306), .B0(n1046), .B1(n303), .C0(n479), 
        .Y(n645) );
  OA22X1 U1067 ( .A0(n333), .A1(n1140), .B0(n302), .B1(n682), .Y(n479) );
  OAI221XL U1068 ( .A0(n1094), .A1(n306), .B0(n1059), .B1(n303), .C0(n482), 
        .Y(n646) );
  AOI2BB2XL U1069 ( .B0(n319), .B1(MEMWriteData[15]), .A0N(n302), .A1N(n1156), 
        .Y(n482) );
  OAI221XL U1070 ( .A0(n1095), .A1(n306), .B0(n1060), .B1(n303), .C0(n485), 
        .Y(n647) );
  AOI2BB2XL U1071 ( .B0(n319), .B1(MEMWriteData[14]), .A0N(n302), .A1N(n1168), 
        .Y(n485) );
  OAI221XL U1072 ( .A0(n1096), .A1(n306), .B0(n1061), .B1(n303), .C0(n488), 
        .Y(n648) );
  AOI2BB2XL U1073 ( .B0(n319), .B1(MEMWriteData[13]), .A0N(n302), .A1N(n1162), 
        .Y(n488) );
  OAI221XL U1074 ( .A0(n1097), .A1(n306), .B0(n1062), .B1(n303), .C0(n491), 
        .Y(n649) );
  AOI2BB2XL U1075 ( .B0(n319), .B1(MEMWriteData[12]), .A0N(n302), .A1N(n1159), 
        .Y(n491) );
  OAI221XL U1076 ( .A0(n1098), .A1(n306), .B0(n1063), .B1(n303), .C0(n494), 
        .Y(n650) );
  AOI2BB2XL U1077 ( .B0(n319), .B1(MEMWriteData[11]), .A0N(n302), .A1N(n1165), 
        .Y(n494) );
  OAI221XL U1078 ( .A0(n1092), .A1(n305), .B0(n1057), .B1(n304), .C0(n527), 
        .Y(n661) );
  AOI2BB2XL U1079 ( .B0(n319), .B1(MEMWriteData[17]), .A0N(n301), .A1N(n693), 
        .Y(n527) );
  OAI221XL U1080 ( .A0(n1091), .A1(n305), .B0(n1056), .B1(n304), .C0(n530), 
        .Y(n662) );
  AOI2BB2XL U1081 ( .B0(n319), .B1(MEMWriteData[18]), .A0N(n301), .A1N(n692), 
        .Y(n530) );
  OAI221XL U1082 ( .A0(n1089), .A1(n305), .B0(n1054), .B1(n304), .C0(n533), 
        .Y(n663) );
  AOI2BB2XL U1083 ( .B0(n319), .B1(MEMWriteData[20]), .A0N(n301), .A1N(n690), 
        .Y(n533) );
  OAI221XL U1084 ( .A0(n1080), .A1(n305), .B0(n1045), .B1(n304), .C0(n536), 
        .Y(n664) );
  OA22X1 U1085 ( .A0(n332), .A1(n1137), .B0(n302), .B1(n681), .Y(n536) );
  OAI221XL U1086 ( .A0(n1093), .A1(n305), .B0(n1058), .B1(n303), .C0(n539), 
        .Y(n665) );
  AOI2BB2XL U1087 ( .B0(n319), .B1(MEMWriteData[16]), .A0N(n301), .A1N(n694), 
        .Y(n539) );
  OAI221XL U1088 ( .A0(n1079), .A1(n305), .B0(n1044), .B1(n304), .C0(n542), 
        .Y(n666) );
  OA22X1 U1089 ( .A0(n333), .A1(n1134), .B0(n301), .B1(n680), .Y(n542) );
  OAI221XL U1090 ( .A0(n1078), .A1(n305), .B0(n1043), .B1(n303), .C0(n545), 
        .Y(n667) );
  OA22X1 U1091 ( .A0(n332), .A1(n1130), .B0(n301), .B1(n679), .Y(n545) );
  OAI221XL U1092 ( .A0(n1099), .A1(n306), .B0(n1064), .B1(n303), .C0(n497), 
        .Y(n651) );
  AOI2BB2XL U1093 ( .B0(n319), .B1(MEMWriteData[10]), .A0N(n302), .A1N(n1180), 
        .Y(n497) );
  OAI221XL U1094 ( .A0(n1100), .A1(n306), .B0(n1065), .B1(n303), .C0(n500), 
        .Y(n652) );
  AOI2BB2XL U1095 ( .B0(n319), .B1(MEMWriteData[9]), .A0N(n301), .A1N(n1171), 
        .Y(n500) );
  OAI221XL U1096 ( .A0(n1101), .A1(n306), .B0(n1066), .B1(n303), .C0(n503), 
        .Y(n653) );
  AOI2BB2XL U1097 ( .B0(n319), .B1(MEMWriteData[8]), .A0N(n301), .A1N(n703), 
        .Y(n503) );
  OAI221XL U1098 ( .A0(n1102), .A1(n305), .B0(n1067), .B1(n303), .C0(n506), 
        .Y(n654) );
  AOI2BB2XL U1099 ( .B0(n319), .B1(MEMWriteData[7]), .A0N(n301), .A1N(n1174), 
        .Y(n506) );
  OAI221XL U1100 ( .A0(n1103), .A1(n305), .B0(n1068), .B1(n304), .C0(n509), 
        .Y(n655) );
  AOI2BB2XL U1101 ( .B0(n319), .B1(MEMWriteData[6]), .A0N(n301), .A1N(n1186), 
        .Y(n509) );
  OAI221XL U1102 ( .A0(n1104), .A1(n305), .B0(n1069), .B1(n303), .C0(n512), 
        .Y(n656) );
  AOI2BB2XL U1103 ( .B0(n321), .B1(MEMWriteData[5]), .A0N(n301), .A1N(n1177), 
        .Y(n512) );
  OAI221XL U1104 ( .A0(n1105), .A1(n305), .B0(n1070), .B1(n304), .C0(n515), 
        .Y(n657) );
  AOI2BB2XL U1105 ( .B0(n320), .B1(MEMWriteData[4]), .A0N(n301), .A1N(n842), 
        .Y(n515) );
  OAI221XL U1106 ( .A0(n1106), .A1(n305), .B0(n1071), .B1(n453), .C0(n518), 
        .Y(n658) );
  AOI2BB2XL U1107 ( .B0(n319), .B1(MEMWriteData[3]), .A0N(n301), .A1N(n1153), 
        .Y(n518) );
  OAI221XL U1108 ( .A0(n1107), .A1(n305), .B0(n1072), .B1(n303), .C0(n521), 
        .Y(n659) );
  AOI2BB2XL U1109 ( .B0(n320), .B1(MEMWriteData[2]), .A0N(n301), .A1N(n1183), 
        .Y(n521) );
  NOR2BX1 U1110 ( .AN(n332), .B(ID_EX[4]), .Y(n162) );
  AND2X2 U1111 ( .A(ID_EX[4]), .B(n332), .Y(n163) );
  OAI2BB2XL U1112 ( .B0(n632), .B1(n333), .A0N(ID_MEM[0]), .A1N(n333), .Y(n669) );
  OAI2BB2XL U1113 ( .B0(n633), .B1(n333), .A0N(ID_MEM[1]), .A1N(n333), .Y(n670) );
  OAI2BB2XL U1114 ( .B0(n634), .B1(n333), .A0N(ID_MEM[2]), .A1N(n333), .Y(n671) );
  OAI2BB2XL U1115 ( .B0(n635), .B1(n333), .A0N(ID_WB[0]), .A1N(n333), .Y(n672)
         );
  CLKMX2X2 U1116 ( .A(ID_WB[1]), .B(n1146), .S0(n320), .Y(n673) );
  OAI221X2 U1117 ( .A0(n679), .A1(n277), .B0(n1043), .B1(n273), .C0(n363), .Y(
        ALUData1[31]) );
  OAI221X2 U1118 ( .A0(n680), .A1(n277), .B0(n1044), .B1(n273), .C0(n365), .Y(
        ALUData1[30]) );
  OAI221X2 U1119 ( .A0(n681), .A1(n277), .B0(n1045), .B1(n273), .C0(n366), .Y(
        ALUData1[29]) );
  OAI221X2 U1120 ( .A0(n682), .A1(n277), .B0(n1046), .B1(n273), .C0(n369), .Y(
        ALUData1[28]) );
  OAI221X2 U1121 ( .A0(n683), .A1(n277), .B0(n1047), .B1(n273), .C0(n370), .Y(
        ALUData1[27]) );
  NAND3BX2 U1122 ( .AN(n372), .B(n444), .C(n1042), .Y(n1013) );
  OAI221X2 U1123 ( .A0(n684), .A1(n277), .B0(n1048), .B1(n273), .C0(n394), .Y(
        ALUData1[26]) );
  OAI221X2 U1124 ( .A0(n685), .A1(n277), .B0(n1049), .B1(n273), .C0(n409), .Y(
        ALUData1[25]) );
  OAI221X2 U1125 ( .A0(n686), .A1(n277), .B0(n1050), .B1(n273), .C0(n426), .Y(
        ALUData1[24]) );
  OAI221X2 U1126 ( .A0(n687), .A1(n277), .B0(n1051), .B1(n273), .C0(n466), .Y(
        ALUData1[23]) );
  OAI221X2 U1127 ( .A0(n688), .A1(n277), .B0(n1052), .B1(n273), .C0(n493), .Y(
        ALUData1[22]) );
  OAI221X2 U1128 ( .A0(n689), .A1(n277), .B0(n1053), .B1(n273), .C0(n522), .Y(
        ALUData1[21]) );
  OAI221X2 U1129 ( .A0(n690), .A1(n277), .B0(n1054), .B1(n273), .C0(n552), .Y(
        ALUData1[20]) );
  OAI221X2 U1130 ( .A0(n691), .A1(n277), .B0(n1055), .B1(n273), .C0(n570), .Y(
        ALUData1[19]) );
  CLKINVX3 U1131 ( .A(n251), .Y(n1018) );
  OAI221X2 U1132 ( .A0(n692), .A1(n276), .B0(n1056), .B1(n273), .C0(n591), .Y(
        ALUData1[18]) );
  OAI221X2 U1133 ( .A0(n693), .A1(n275), .B0(n1057), .B1(n273), .C0(n615), .Y(
        ALUData1[17]) );
  OAI221X2 U1134 ( .A0(n694), .A1(n276), .B0(n1058), .B1(n273), .C0(n719), .Y(
        ALUData1[16]) );
  OAI221X2 U1135 ( .A0(n1157), .A1(n275), .B0(n1059), .B1(n273), .C0(n747), 
        .Y(ALUData1[15]) );
  OAI221X2 U1136 ( .A0(n1169), .A1(n276), .B0(n1060), .B1(n273), .C0(n749), 
        .Y(ALUData1[14]) );
  OAI221X2 U1137 ( .A0(n1163), .A1(n276), .B0(n1061), .B1(n273), .C0(n762), 
        .Y(ALUData1[13]) );
  OAI221X2 U1138 ( .A0(n1160), .A1(n275), .B0(n1062), .B1(n273), .C0(n775), 
        .Y(ALUData1[12]) );
  OAI221X2 U1139 ( .A0(n1166), .A1(n275), .B0(n1063), .B1(n273), .C0(n788), 
        .Y(ALUData1[11]) );
  OAI221X2 U1140 ( .A0(n1180), .A1(n276), .B0(n1064), .B1(n273), .C0(n802), 
        .Y(ALUData1[10]) );
  OAI221X2 U1141 ( .A0(n1172), .A1(n275), .B0(n1065), .B1(n273), .C0(n815), 
        .Y(n702) );
  OAI221X2 U1142 ( .A0(n703), .A1(n275), .B0(n1066), .B1(n273), .C0(n828), .Y(
        ALUData1[8]) );
  OAI221X2 U1143 ( .A0(n1174), .A1(n276), .B0(n1067), .B1(n274), .C0(n840), 
        .Y(ALUData1[7]) );
  OAI221X2 U1144 ( .A0(n1186), .A1(n275), .B0(n1068), .B1(n274), .C0(n853), 
        .Y(ALUData1[6]) );
  OAI221X2 U1145 ( .A0(n1177), .A1(n276), .B0(n1069), .B1(n274), .C0(n865), 
        .Y(ALUData1[5]) );
  OAI221X2 U1146 ( .A0(n855), .A1(n276), .B0(n1070), .B1(n274), .C0(n878), .Y(
        ALUData1[4]) );
  OAI221X2 U1147 ( .A0(n842), .A1(n283), .B0(n250), .B1(n1116), .C0(n879), .Y(
        ALUData2[4]) );
  OAI221X2 U1148 ( .A0(n1184), .A1(n276), .B0(n1072), .B1(n274), .C0(n903), 
        .Y(ALUData1[2]) );
  OAI221X2 U1149 ( .A0(n710), .A1(n276), .B0(n274), .B1(n1039), .C0(n915), .Y(
        ALUData1[1]) );
  OAI221X2 U1150 ( .A0(n1149), .A1(n276), .B0(n274), .B1(n1035), .C0(n929), 
        .Y(ALUData1[0]) );
  Execution_DW_cmp_0 lte_117 ( .A({ALUData1[31:10], n702, ALUData1[8:0]}), .B(
        {n251, n252, n253, n254, n255, n259, n260, n261, n262, n263, n264, 
        n265, n266, n267, n270, n271, ALUData2[15], n108, ALUData2[13:12], 
        n134, ALUData2[10:1], n5}), .TC(1'b0), .GE_LT(1'b0), .GE_GT_EQ(1'b0), 
        .GE_LT_GT_LE(N524) );
  Execution_DW_rightsh_0 srl_80 ( .A({n251, n252, n253, n254, n255, n259, n260, 
        n261, n262, n263, n264, n265, n266, n267, n270, n271, ALUData2[15], 
        n108, ALUData2[13:12], n134, ALUData2[10:1], n5}), .DATA_TC(1'b0), 
        .SH({n317, n315, n311, n309, n307}), .B({N395, N394, N393, N392, N391, 
        N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, 
        N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, 
        N366, N365, N364}) );
  Execution_DW_leftsh_0 sll_79 ( .A({n251, n252, n253, n254, n255, n259, n260, 
        n261, n262, n263, n264, n265, n266, n267, n270, n271, ALUData2[15], 
        n108, ALUData2[13:12], n134, ALUData2[10:1], n5}), .SH({n317, n315, 
        n311, n309, n307}), .B({N363, N362, N361, N360, N359, N358, N357, N356, 
        N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344, 
        N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, N332}) );
  Execution_DW01_sub_1 sub_74 ( .A({ALUData1[31:10], n702, ALUData1[8:0]}), 
        .B({n251, n252, n253, n254, n255, n259, n260, n261, n262, n263, n264, 
        n265, n266, n267, n270, n271, ALUData2[15], n108, ALUData2[13:1], n5}), 
        .CI(1'b0), .DIFF({N235, N234, N233, N232, N231, N230, N229, N228, N227, 
        N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, 
        N214, N213, N212, N211, N210, N209, N208, N207, N206, N205, N204}) );
  Execution_DW01_add_1 add_73 ( .A({ALUData1[31:10], n702, ALUData1[8:0]}), 
        .B({n251, n252, n253, n254, n255, n259, n260, n261, n262, n263, n264, 
        n265, n266, n267, n270, n271, ALUData2[15], n108, ALUData2[13:1], n5}), 
        .CI(1'b0), .SUM({N203, N202, N201, N200, N199, N198, N197, N196, N195, 
        N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, 
        N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172}) );
  INVXL U160 ( .A(n1131), .Y(n1129) );
  INVX12 U1151 ( .A(n1129), .Y(MEMWriteData[1]) );
  SDFFRXL \WB_reg[0]  ( .D(n672), .SI(n36), .SE(test_se), .CK(clk), .RN(n345), 
        .Q(WB[0]), .QN(n635) );
  SDFFRXL \MEM_reg[2]  ( .D(n671), .SI(n633), .SE(test_se), .CK(clk), .RN(n345), .Q(MEM[2]), .QN(n634) );
  SDFFRXL \ALUresult_reg[14]  ( .D(next_ALUresult[14]), .SI(n90), .SE(test_se), 
        .CK(clk), .RN(n341), .Q(n92), .QN(n696) );
  SDFFRXL \ALUresult_reg[11]  ( .D(next_ALUresult[11]), .SI(n86), .SE(test_se), 
        .CK(clk), .RN(n342), .Q(n91), .QN(n699) );
  SDFFRXL \ALUresult_reg[13]  ( .D(next_ALUresult[13]), .SI(n84), .SE(test_se), 
        .CK(clk), .RN(n341), .Q(n90), .QN(n697) );
  SDFFRXL \ALUresult_reg[6]  ( .D(next_ALUresult[6]), .SI(n85), .SE(test_se), 
        .CK(clk), .RN(n343), .Q(n89), .QN(n705) );
  SDFFRXL \ALUresult_reg[3]  ( .D(next_ALUresult[3]), .SI(n87), .SE(test_se), 
        .CK(clk), .RN(n343), .Q(n88), .QN(n708) );
  SDFFRXL \ALUresult_reg[2]  ( .D(next_ALUresult[2]), .SI(ALUresult[1]), .SE(
        test_se), .CK(clk), .RN(n343), .Q(n87), .QN(n709) );
  SDFFRXL \ALUresult_reg[10]  ( .D(next_ALUresult[10]), .SI(n81), .SE(test_se), 
        .CK(clk), .RN(n342), .Q(n86), .QN(n700) );
  SDFFRXL \ALUresult_reg[24]  ( .D(next_ALUresult[24]), .SI(ALUresult[23]), 
        .SE(test_se), .CK(clk), .RN(n340), .Q(n430), .QN(n686) );
  SDFFRXL \ALUresult_reg[27]  ( .D(next_ALUresult[27]), .SI(ALUresult[26]), 
        .SE(test_se), .CK(clk), .RN(n341), .Q(n1122), .QN(n683) );
  SDFFRXL \ALUresult_reg[22]  ( .D(next_ALUresult[22]), .SI(ALUresult[21]), 
        .SE(test_se), .CK(clk), .RN(n340), .Q(n1125), .QN(n688) );
  SDFFRXL \ALUresult_reg[5]  ( .D(next_ALUresult[5]), .SI(ALUresult[4]), .SE(
        test_se), .CK(clk), .RN(n343), .Q(n85), .QN(n706) );
  SDFFRXL \ALUresult_reg[25]  ( .D(next_ALUresult[25]), .SI(ALUresult[24]), 
        .SE(test_se), .CK(clk), .RN(n340), .Q(n411), .QN(n685) );
  SDFFRXL \ALUresult_reg[31]  ( .D(next_ALUresult[31]), .SI(ALUresult[30]), 
        .SE(test_se), .CK(clk), .RN(n345), .Q(n1121), .QN(n679) );
  SDFFRXL \ALUresult_reg[26]  ( .D(next_ALUresult[26]), .SI(ALUresult[25]), 
        .SE(test_se), .CK(clk), .RN(n341), .Q(n1123), .QN(n684) );
  SDFFRXL \ALUresult_reg[23]  ( .D(next_ALUresult[23]), .SI(ALUresult[22]), 
        .SE(test_se), .CK(clk), .RN(n340), .Q(n1124), .QN(n687) );
  SDFFRXL \ALUresult_reg[18]  ( .D(next_ALUresult[18]), .SI(ALUresult[17]), 
        .SE(test_se), .CK(clk), .RN(n344), .Q(n1127), .QN(n692) );
  SDFFRXL \ALUresult_reg[19]  ( .D(next_ALUresult[19]), .SI(ALUresult[18]), 
        .SE(test_se), .CK(clk), .RN(n340), .Q(n1126), .QN(n691) );
  SDFFRXL \ALUresult_reg[12]  ( .D(next_ALUresult[12]), .SI(n91), .SE(test_se), 
        .CK(clk), .RN(n342), .Q(n84), .QN(n698) );
  SDFFRXL \ALUresult_reg[7]  ( .D(next_ALUresult[7]), .SI(n89), .SE(test_se), 
        .CK(clk), .RN(n342), .Q(n83), .QN(n704) );
  SDFFRXL \ALUresult_reg[15]  ( .D(next_ALUresult[15]), .SI(n92), .SE(test_se), 
        .CK(clk), .RN(n341), .Q(n82), .QN(n695) );
  SDFFRXL \ALUresult_reg[9]  ( .D(next_ALUresult[9]), .SI(ALUresult[8]), .SE(
        test_se), .CK(clk), .RN(n342), .Q(n81), .QN(n701) );
  SDFFRXL \ALUresult_reg[0]  ( .D(next_ALUresult[0]), .SI(test_si), .SE(
        test_se), .CK(clk), .RN(n345), .Q(n1128), .QN(n711) );
  SDFFRXL \MEM_reg[1]  ( .D(n670), .SI(n632), .SE(test_se), .CK(clk), .RN(n345), .Q(MEM[1]), .QN(n633) );
  SDFFRXL \MEM_reg[0]  ( .D(n669), .SI(n41), .SE(test_se), .CK(clk), .RN(n345), 
        .Q(MEM[0]), .QN(n632) );
  SDFFRXL \MEMWriteData_reg[19]  ( .D(n637), .SI(n48), .SE(test_se), .CK(clk), 
        .RN(n340), .Q(n80), .QN(n11) );
  SDFFRXL \MEMWriteData_reg[21]  ( .D(n638), .SI(n47), .SE(test_se), .CK(clk), 
        .RN(n340), .Q(n78), .QN(n12) );
  SDFFRXL \MEMWriteData_reg[22]  ( .D(n639), .SI(n78), .SE(test_se), .CK(clk), 
        .RN(n340), .Q(n76), .QN(n13) );
  SDFFRXL \MEMWriteData_reg[23]  ( .D(n640), .SI(n76), .SE(test_se), .CK(clk), 
        .RN(n340), .Q(n74), .QN(n14) );
  SDFFRXL \MEMWriteData_reg[24]  ( .D(n641), .SI(n74), .SE(test_se), .CK(clk), 
        .RN(n340), .Q(n72), .QN(n15) );
  SDFFRXL \MEMWriteData_reg[25]  ( .D(n642), .SI(n72), .SE(test_se), .CK(clk), 
        .RN(n340), .Q(n70), .QN(n16) );
  SDFFRXL \MEMWriteData_reg[26]  ( .D(n643), .SI(n70), .SE(test_se), .CK(clk), 
        .RN(n341), .Q(n68), .QN(n17) );
  SDFFRXL \MEMWriteData_reg[15]  ( .D(n646), .SI(n64), .SE(test_se), .CK(clk), 
        .RN(n341), .Q(n66), .QN(n18) );
  SDFFRXL \MEMWriteData_reg[14]  ( .D(n647), .SI(n62), .SE(test_se), .CK(clk), 
        .RN(n341), .Q(n64), .QN(n19) );
  SDFFRXL \MEMWriteData_reg[13]  ( .D(n648), .SI(n60), .SE(test_se), .CK(clk), 
        .RN(n341), .Q(n62), .QN(n20) );
  SDFFRXL \MEMWriteData_reg[12]  ( .D(n649), .SI(n59), .SE(test_se), .CK(clk), 
        .RN(n342), .Q(n60), .QN(n21) );
  SDFFRXL \MEMWriteData_reg[11]  ( .D(n650), .SI(n58), .SE(test_se), .CK(clk), 
        .RN(n342), .Q(n59), .QN(n22) );
  SDFFRXL \MEMWriteData_reg[10]  ( .D(n651), .SI(n57), .SE(test_se), .CK(clk), 
        .RN(n342), .Q(n58), .QN(n27) );
  SDFFRXL \MEMWriteData_reg[9]  ( .D(n652), .SI(n56), .SE(test_se), .CK(clk), 
        .RN(n342), .Q(n57), .QN(n28) );
  SDFFRXL \MEMWriteData_reg[8]  ( .D(n653), .SI(n55), .SE(test_se), .CK(clk), 
        .RN(n342), .Q(n56), .QN(n29) );
  SDFFRXL \MEMWriteData_reg[7]  ( .D(n654), .SI(n54), .SE(test_se), .CK(clk), 
        .RN(n342), .Q(n55), .QN(n30) );
  SDFFRXL \MEMWriteData_reg[6]  ( .D(n655), .SI(n53), .SE(test_se), .CK(clk), 
        .RN(n343), .Q(n54), .QN(n31) );
  SDFFRXL \MEMWriteData_reg[5]  ( .D(n656), .SI(n52), .SE(test_se), .CK(clk), 
        .RN(n343), .Q(n53), .QN(n32) );
  SDFFRXL \MEMWriteData_reg[4]  ( .D(n657), .SI(n51), .SE(test_se), .CK(clk), 
        .RN(n343), .Q(n52), .QN(n33) );
  SDFFRXL \MEMWriteData_reg[3]  ( .D(n658), .SI(n50), .SE(test_se), .CK(clk), 
        .RN(n343), .Q(n51), .QN(n34) );
  SDFFRXL \MEMWriteData_reg[2]  ( .D(n659), .SI(n1037), .SE(test_se), .CK(clk), 
        .RN(n343), .Q(n50), .QN(n35) );
  SDFFRXL \MEMWriteData_reg[17]  ( .D(n661), .SI(n46), .SE(test_se), .CK(clk), 
        .RN(n344), .Q(n49), .QN(n23) );
  SDFFRXL \MEMWriteData_reg[18]  ( .D(n662), .SI(n49), .SE(test_se), .CK(clk), 
        .RN(n344), .Q(n48), .QN(n24) );
  SDFFRXL \MEMWriteData_reg[20]  ( .D(n663), .SI(n80), .SE(test_se), .CK(clk), 
        .RN(n344), .Q(n47), .QN(n25) );
  SDFFRXL \MEMWriteData_reg[16]  ( .D(n665), .SI(n66), .SE(test_se), .CK(clk), 
        .RN(n344), .Q(n46), .QN(n26) );
  SDFFRXL \MEMWriteData_reg[27]  ( .D(n644), .SI(n68), .SE(test_se), .CK(clk), 
        .RN(n341), .Q(n45), .QN(n1031) );
  SDFFRXL \MEMWriteData_reg[28]  ( .D(n645), .SI(n45), .SE(test_se), .CK(clk), 
        .RN(n341), .Q(n44), .QN(n1030) );
  SDFFRXL \MEMWriteData_reg[29]  ( .D(n664), .SI(n44), .SE(test_se), .CK(clk), 
        .RN(n344), .Q(n43), .QN(n1029) );
  SDFFRXL \MEMWriteData_reg[30]  ( .D(n666), .SI(n43), .SE(test_se), .CK(clk), 
        .RN(n344), .Q(n42), .QN(n1028) );
  SDFFRXL \MEMWriteData_reg[31]  ( .D(n667), .SI(n42), .SE(test_se), .CK(clk), 
        .RN(n345), .Q(n41), .QN(n1027) );
  SDFFRXL \MEMWriteData_reg[0]  ( .D(n668), .SI(ALUresult[31]), .SE(test_se), 
        .CK(clk), .RN(n345), .Q(n40), .QN(n1033) );
  SDFFRXL \RegisterRd_reg[2]  ( .D(n1075), .SI(n3), .SE(test_se), .CK(clk), 
        .RN(rst), .Q(n1191), .QN(n39) );
  SDFFRXL \RegisterRd_reg[0]  ( .D(n1077), .SI(MEM[2]), .SE(test_se), .CK(clk), 
        .RN(n345), .Q(n1192), .QN(n38) );
  SDFFRXL \ALUresult_reg[1]  ( .D(next_ALUresult[1]), .SI(ALUresult[0]), .SE(
        test_se), .CK(clk), .RN(n343), .Q(n917), .QN(n710) );
  SDFFRXL \ALUresult_reg[8]  ( .D(next_ALUresult[8]), .SI(n83), .SE(test_se), 
        .CK(clk), .RN(n342), .Q(n829), .QN(n703) );
  SDFFRXL \ALUresult_reg[21]  ( .D(next_ALUresult[21]), .SI(ALUresult[20]), 
        .SE(test_se), .CK(clk), .RN(n340), .Q(n524), .QN(n689) );
  SDFFRXL \ALUresult_reg[20]  ( .D(next_ALUresult[20]), .SI(ALUresult[19]), 
        .SE(test_se), .CK(clk), .RN(n344), .Q(n554), .QN(n690) );
  SDFFRXL \ALUresult_reg[28]  ( .D(next_ALUresult[28]), .SI(ALUresult[27]), 
        .SE(test_se), .CK(clk), .RN(n341), .Q(n961), .QN(n682) );
  SDFFRXL \ALUresult_reg[29]  ( .D(next_ALUresult[29]), .SI(ALUresult[28]), 
        .SE(test_se), .CK(clk), .RN(n344), .Q(n974), .QN(n681) );
  SDFFRXL \ALUresult_reg[16]  ( .D(next_ALUresult[16]), .SI(n82), .SE(test_se), 
        .CK(clk), .RN(n344), .Q(n721), .QN(n694) );
  SDFFRXL \ALUresult_reg[4]  ( .D(next_ALUresult[4]), .SI(n88), .SE(test_se), 
        .CK(clk), .RN(n343), .Q(n880), .QN(n707) );
  SDFFRXL \ALUresult_reg[17]  ( .D(next_ALUresult[17]), .SI(ALUresult[16]), 
        .SE(test_se), .CK(clk), .RN(n344), .Q(n617), .QN(n693) );
  SDFFRXL \ALUresult_reg[30]  ( .D(next_ALUresult[30]), .SI(ALUresult[29]), 
        .SE(test_se), .CK(clk), .RN(n344), .Q(n990), .QN(n680) );
  SDFFRXL \WB_reg[1]  ( .D(n673), .SI(n635), .SE(test_se), .CK(clk), .RN(n345), 
        .Q(n1189), .QN(test_so) );
  SDFFRXL \RegisterRd_reg[4]  ( .D(n1073), .SI(n4), .SE(test_se), .CK(clk), 
        .RN(n346), .Q(n1190), .QN(n36) );
  SDFFRX2 \RegisterRd_reg[3]  ( .D(n1074), .SI(n39), .SE(test_se), .CK(clk), 
        .RN(n346), .Q(RegisterRd[3]), .QN(n4) );
  SDFFRX2 \RegisterRd_reg[1]  ( .D(n1076), .SI(n38), .SE(test_se), .CK(clk), 
        .RN(n345), .Q(RegisterRd[1]), .QN(n3) );
  SDFFRXL \MEMWriteData_reg[1]  ( .D(n660), .SI(n40), .SE(test_se), .CK(clk), 
        .RN(rst), .Q(n1131), .QN(n1037) );
  CLKBUFX2 U1 ( .A(n708), .Y(n93) );
  CLKBUFX2 U2 ( .A(n695), .Y(n94) );
  CLKBUFX2 U7 ( .A(n698), .Y(n95) );
  CLKBUFX2 U8 ( .A(n697), .Y(n96) );
  CLKBUFX2 U9 ( .A(n699), .Y(n97) );
  CLKBUFX2 U10 ( .A(n696), .Y(n98) );
  CLKBUFX2 U1152 ( .A(n701), .Y(n104) );
  CLKBUFX2 U1153 ( .A(n704), .Y(n751) );
  CLKBUFX2 U1154 ( .A(n706), .Y(n764) );
  CLKBUFX2 U1155 ( .A(n700), .Y(n777) );
  CLKBUFX2 U1156 ( .A(n709), .Y(n791) );
  CLKBUFX2 U1157 ( .A(n705), .Y(n804) );
  INVXL U1158 ( .A(n707), .Y(n817) );
  INVXL U1159 ( .A(n817), .Y(n842) );
  INVXL U1160 ( .A(n817), .Y(n855) );
  INVXL U1161 ( .A(n1033), .Y(n868) );
  INVXL U1162 ( .A(n868), .Y(n892) );
  INVXL U1163 ( .A(n868), .Y(n905) );
  INVXL U1164 ( .A(n1027), .Y(n950) );
  INVXL U1165 ( .A(n950), .Y(n1041) );
  INVXL U1166 ( .A(n950), .Y(n1130) );
  INVXL U1167 ( .A(n1028), .Y(n1132) );
  INVXL U1168 ( .A(n1132), .Y(n1133) );
  INVXL U1169 ( .A(n1132), .Y(n1134) );
  INVXL U1170 ( .A(n1029), .Y(n1135) );
  INVXL U1171 ( .A(n1135), .Y(n1136) );
  INVXL U1172 ( .A(n1135), .Y(n1137) );
  INVXL U1173 ( .A(n1030), .Y(n1138) );
  INVXL U1174 ( .A(n1138), .Y(n1139) );
  INVXL U1175 ( .A(n1138), .Y(n1140) );
  INVXL U1176 ( .A(n1031), .Y(n1141) );
  INVXL U1177 ( .A(n1141), .Y(n1142) );
  INVXL U1178 ( .A(n1141), .Y(n1143) );
  INVXL U1179 ( .A(n1189), .Y(n1144) );
  INVXL U1180 ( .A(n1144), .Y(WB[1]) );
  INVXL U1181 ( .A(n1144), .Y(n1146) );
  INVXL U1182 ( .A(n711), .Y(n1147) );
  INVXL U1183 ( .A(n1147), .Y(n1148) );
  INVXL U1184 ( .A(n1147), .Y(n1149) );
  CLKBUFX2 U1185 ( .A(n1191), .Y(RegisterRd[2]) );
  CLKBUFX2 U1186 ( .A(n1192), .Y(RegisterRd[0]) );
  INVXL U1187 ( .A(n708), .Y(n1152) );
  INVXL U1188 ( .A(n1152), .Y(n1153) );
  INVXL U1189 ( .A(n1152), .Y(n1154) );
  INVXL U1190 ( .A(n695), .Y(n1155) );
  INVXL U1191 ( .A(n1155), .Y(n1156) );
  INVXL U1192 ( .A(n1155), .Y(n1157) );
  INVXL U1193 ( .A(n698), .Y(n1158) );
  INVXL U1194 ( .A(n1158), .Y(n1159) );
  INVXL U1195 ( .A(n1158), .Y(n1160) );
  INVXL U1196 ( .A(n697), .Y(n1161) );
  INVXL U1197 ( .A(n1161), .Y(n1162) );
  INVXL U1198 ( .A(n1161), .Y(n1163) );
  INVXL U1199 ( .A(n699), .Y(n1164) );
  INVXL U1200 ( .A(n1164), .Y(n1165) );
  INVXL U1201 ( .A(n1164), .Y(n1166) );
  INVXL U1202 ( .A(n696), .Y(n1167) );
  INVXL U1203 ( .A(n1167), .Y(n1168) );
  INVXL U1204 ( .A(n1167), .Y(n1169) );
  INVXL U1205 ( .A(n701), .Y(n1170) );
  INVXL U1206 ( .A(n1170), .Y(n1171) );
  INVXL U1207 ( .A(n1170), .Y(n1172) );
  INVXL U1208 ( .A(n704), .Y(n1173) );
  INVXL U1209 ( .A(n1173), .Y(n1174) );
  INVXL U1210 ( .A(n1173), .Y(n1175) );
  INVXL U1211 ( .A(n706), .Y(n1176) );
  INVXL U1212 ( .A(n1176), .Y(n1177) );
  INVXL U1213 ( .A(n1176), .Y(n1178) );
  INVXL U1214 ( .A(n700), .Y(n1179) );
  INVXL U1215 ( .A(n1179), .Y(n1180) );
  INVXL U1216 ( .A(n1179), .Y(n1181) );
  INVXL U1217 ( .A(n709), .Y(n1182) );
  INVXL U1218 ( .A(n1182), .Y(n1183) );
  INVXL U1219 ( .A(n1182), .Y(n1184) );
  INVXL U1220 ( .A(n705), .Y(n1185) );
  INVXL U1221 ( .A(n1185), .Y(n1186) );
  INVXL U1222 ( .A(n1185), .Y(n1187) );
  CLKBUFX2 U1223 ( .A(n1190), .Y(RegisterRd[4]) );
endmodule


module InstructionDecode_DW_mult_uns_1 ( a, b, product );
  input [31:0] a;
  output [32:0] product;
  input b;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33;

  CLKBUFX12 U67 ( .A(n33), .Y(n2) );
  NOR2X2 U68 ( .A(n1), .B(n20), .Y(product[14]) );
  NOR2X1 U69 ( .A(n2), .B(n17), .Y(product[17]) );
  NOR2X1 U70 ( .A(n1), .B(n24), .Y(product[10]) );
  NOR2X1 U71 ( .A(n1), .B(n18), .Y(product[16]) );
  NOR2X1 U72 ( .A(n2), .B(n11), .Y(product[23]) );
  NOR2X1 U73 ( .A(n1), .B(n21), .Y(product[13]) );
  NOR2X1 U74 ( .A(n2), .B(n15), .Y(product[19]) );
  NOR2X1 U75 ( .A(n1), .B(n25), .Y(product[9]) );
  NOR2X1 U76 ( .A(n2), .B(n9), .Y(product[25]) );
  NOR2X1 U77 ( .A(n2), .B(n10), .Y(product[24]) );
  NOR2X1 U78 ( .A(n1), .B(n22), .Y(product[12]) );
  NOR2X1 U79 ( .A(n1), .B(n27), .Y(product[7]) );
  NOR2X1 U80 ( .A(n1), .B(n32), .Y(product[2]) );
  NOR2X1 U81 ( .A(n1), .B(n26), .Y(product[8]) );
  NOR2X1 U82 ( .A(n1), .B(n28), .Y(product[6]) );
  CLKINVX4 U83 ( .A(b), .Y(n33) );
  NOR2X1 U84 ( .A(n2), .B(n12), .Y(product[22]) );
  BUFX12 U85 ( .A(n33), .Y(n1) );
  NOR2XL U86 ( .A(n1), .B(n30), .Y(product[4]) );
  NOR2XL U87 ( .A(n2), .B(n14), .Y(product[20]) );
  NOR2XL U88 ( .A(n2), .B(n13), .Y(product[21]) );
  NOR2XL U89 ( .A(n1), .B(n29), .Y(product[5]) );
  NOR2XL U90 ( .A(n2), .B(n8), .Y(product[26]) );
  NOR2XL U91 ( .A(n2), .B(n7), .Y(product[27]) );
  NOR2XL U92 ( .A(n2), .B(n6), .Y(product[28]) );
  NOR2XL U93 ( .A(n2), .B(n5), .Y(product[29]) );
  NOR2XL U94 ( .A(n2), .B(n4), .Y(product[30]) );
  NOR2XL U95 ( .A(n2), .B(n3), .Y(product[31]) );
  CLKINVX1 U96 ( .A(a[5]), .Y(n29) );
  CLKINVX1 U97 ( .A(a[7]), .Y(n27) );
  CLKINVX1 U98 ( .A(a[9]), .Y(n25) );
  CLKINVX1 U99 ( .A(a[17]), .Y(n17) );
  NOR2X1 U100 ( .A(n1), .B(n19), .Y(product[15]) );
  CLKINVX1 U101 ( .A(a[15]), .Y(n19) );
  CLKINVX1 U102 ( .A(a[13]), .Y(n21) );
  NOR2X1 U103 ( .A(n1), .B(n23), .Y(product[11]) );
  CLKINVX1 U104 ( .A(a[11]), .Y(n23) );
  CLKINVX1 U105 ( .A(a[23]), .Y(n11) );
  CLKINVX1 U106 ( .A(a[21]), .Y(n13) );
  CLKINVX1 U107 ( .A(a[19]), .Y(n15) );
  CLKINVX1 U108 ( .A(a[27]), .Y(n7) );
  CLKINVX1 U109 ( .A(a[29]), .Y(n5) );
  CLKINVX1 U110 ( .A(a[28]), .Y(n6) );
  CLKINVX1 U111 ( .A(a[2]), .Y(n32) );
  NOR2X1 U112 ( .A(n1), .B(n31), .Y(product[3]) );
  CLKINVX1 U113 ( .A(a[3]), .Y(n31) );
  CLKINVX1 U114 ( .A(a[6]), .Y(n28) );
  CLKINVX1 U115 ( .A(a[12]), .Y(n22) );
  CLKINVX1 U116 ( .A(a[14]), .Y(n20) );
  CLKINVX1 U117 ( .A(a[16]), .Y(n18) );
  NOR2X1 U118 ( .A(n2), .B(n16), .Y(product[18]) );
  CLKINVX1 U119 ( .A(a[18]), .Y(n16) );
  CLKINVX1 U120 ( .A(a[22]), .Y(n12) );
  CLKINVX1 U121 ( .A(a[24]), .Y(n10) );
  CLKINVX1 U122 ( .A(a[25]), .Y(n9) );
  CLKINVX1 U123 ( .A(a[30]), .Y(n4) );
  CLKINVX1 U124 ( .A(a[26]), .Y(n8) );
  CLKINVX1 U125 ( .A(a[4]), .Y(n30) );
  CLKINVX1 U126 ( .A(a[8]), .Y(n26) );
  CLKINVX1 U127 ( .A(a[10]), .Y(n24) );
  CLKINVX1 U128 ( .A(a[20]), .Y(n14) );
  CLKINVX1 U129 ( .A(a[31]), .Y(n3) );
endmodule


module InstructionDecode_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n32, n33, n34, n35, n36, n37, n38, n40, n41, n43, n45, n46, n47, n48,
         n49, n50, n51, n52, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n84, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n116, n117, n118, n119, n120, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n195,
         n196, n197, n198, n199, n201, n202, n203, n205, n207, n209, n212,
         n213, n214, n215, n217, n218, n219, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n348,
         n349, n350, n351, n352, n353, n354, n355, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n1, n31,
         n39, n42, n44, n53, n65, n66, n82, n83, n85, n100, n115, n121;

  NOR2X4 U254 ( .A(n325), .B(A[15]), .Y(n125) );
  NOR2X2 U255 ( .A(n334), .B(A[10]), .Y(n153) );
  BUFX4 U256 ( .A(B[10]), .Y(n334) );
  NOR2X2 U257 ( .A(n86), .B(n59), .Y(n57) );
  BUFX2 U258 ( .A(B[24]), .Y(n321) );
  NOR2X4 U259 ( .A(n118), .B(n113), .Y(n111) );
  NOR2X2 U260 ( .A(B[16]), .B(A[16]), .Y(n118) );
  BUFX4 U261 ( .A(B[11]), .Y(n322) );
  OAI21X2 U262 ( .A0(n125), .A1(n131), .B0(n126), .Y(n124) );
  NOR2X2 U263 ( .A(B[19]), .B(A[19]), .Y(n98) );
  NAND2X2 U264 ( .A(B[6]), .B(A[6]), .Y(n175) );
  OAI21X4 U265 ( .A0(n121), .A1(n184), .B0(n181), .Y(n179) );
  NOR2X8 U267 ( .A(n93), .B(n90), .Y(n88) );
  NOR2X4 U268 ( .A(n332), .B(A[20]), .Y(n93) );
  NAND2X2 U269 ( .A(n334), .B(A[10]), .Y(n154) );
  OAI21X1 U270 ( .A0(n113), .A1(n119), .B0(n114), .Y(n112) );
  OAI21X4 U271 ( .A0(n187), .A1(n190), .B0(n188), .Y(n186) );
  NAND2X2 U272 ( .A(B[2]), .B(A[2]), .Y(n190) );
  CLKBUFX3 U273 ( .A(n176), .Y(n323) );
  NOR2X2 U275 ( .A(n153), .B(n150), .Y(n148) );
  NOR2X4 U276 ( .A(n349), .B(n179), .Y(n177) );
  BUFX8 U277 ( .A(n155), .Y(n324) );
  OAI21X2 U278 ( .A0(n161), .A1(n165), .B0(n162), .Y(n160) );
  NOR2X6 U279 ( .A(n333), .B(n161), .Y(n159) );
  NOR2X2 U280 ( .A(B[9]), .B(A[9]), .Y(n161) );
  NOR2X6 U281 ( .A(n354), .B(n89), .Y(n87) );
  NAND2X4 U282 ( .A(n344), .B(n147), .Y(n145) );
  NAND2X2 U283 ( .A(n342), .B(n343), .Y(n344) );
  CLKINVX1 U284 ( .A(n146), .Y(n343) );
  NOR2X2 U285 ( .A(n324), .B(n134), .Y(n345) );
  XNOR2XL U286 ( .A(n105), .B(n14), .Y(SUM[18]) );
  NAND2X1 U287 ( .A(n123), .B(n111), .Y(n109) );
  AND2X2 U288 ( .A(n186), .B(n178), .Y(n349) );
  NOR2X2 U289 ( .A(n183), .B(n180), .Y(n178) );
  OR2X2 U290 ( .A(n358), .B(n359), .Y(n168) );
  NOR2X1 U291 ( .A(n169), .B(n175), .Y(n358) );
  CLKINVX1 U292 ( .A(n154), .Y(n340) );
  CLKINVX1 U293 ( .A(n324), .Y(n342) );
  CLKBUFX3 U294 ( .A(B[20]), .Y(n332) );
  CLKBUFX3 U295 ( .A(B[21]), .Y(n331) );
  NOR2X1 U296 ( .A(B[22]), .B(A[22]), .Y(n80) );
  NAND2X1 U297 ( .A(n335), .B(A[4]), .Y(n184) );
  CLKBUFX3 U298 ( .A(n164), .Y(n333) );
  AO21X2 U299 ( .A0(n133), .A1(n123), .B0(n124), .Y(n120) );
  NAND2X1 U301 ( .A(B[22]), .B(A[22]), .Y(n81) );
  AO21X1 U303 ( .A0(n145), .A1(n141), .B0(n142), .Y(n363) );
  AOI21X1 U304 ( .A0(n133), .A1(n128), .B0(n129), .Y(n127) );
  XOR2X1 U305 ( .A(n6), .B(n56), .Y(SUM[26]) );
  BUFX4 U306 ( .A(B[15]), .Y(n325) );
  OA21X2 U307 ( .A0(n56), .A1(n54), .B0(n55), .Y(n364) );
  CLKBUFX3 U308 ( .A(B[26]), .Y(n326) );
  OR2X1 U310 ( .A(B[28]), .B(A[28]), .Y(n328) );
  OR2X1 U311 ( .A(B[29]), .B(A[29]), .Y(n329) );
  NOR2X1 U312 ( .A(B[6]), .B(A[6]), .Y(n174) );
  NOR2X1 U313 ( .A(B[14]), .B(A[14]), .Y(n130) );
  CLKINVX1 U314 ( .A(n150), .Y(n339) );
  OAI21X1 U315 ( .A0(n75), .A1(n81), .B0(n76), .Y(n74) );
  NAND2X1 U316 ( .A(B[23]), .B(A[23]), .Y(n76) );
  NAND2X1 U317 ( .A(n330), .B(A[25]), .Y(n64) );
  AOI21X4 U318 ( .A0(n168), .A1(n159), .B0(n160), .Y(n158) );
  NOR2X2 U319 ( .A(n174), .B(n169), .Y(n167) );
  NOR2X2 U320 ( .A(n335), .B(A[4]), .Y(n183) );
  INVXL U321 ( .A(n153), .Y(n212) );
  NOR2X8 U322 ( .A(n355), .B(n108), .Y(n106) );
  OAI21X2 U323 ( .A0(n135), .A1(n109), .B0(n110), .Y(n108) );
  OAI21X2 U324 ( .A0(n90), .A1(n94), .B0(n91), .Y(n89) );
  NOR2X2 U325 ( .A(n331), .B(A[21]), .Y(n90) );
  NAND2XL U326 ( .A(n207), .B(n126), .Y(n17) );
  NAND2X1 U327 ( .A(n325), .B(A[15]), .Y(n126) );
  NOR2X1 U328 ( .A(n348), .B(n112), .Y(n110) );
  INVXL U329 ( .A(n103), .Y(n101) );
  NOR2X4 U330 ( .A(n103), .B(n82), .Y(n96) );
  OAI21X4 U331 ( .A0(n87), .A1(n59), .B0(n60), .Y(n58) );
  AOI21X1 U332 ( .A0(n74), .A1(n61), .B0(n62), .Y(n60) );
  INVX8 U333 ( .A(n106), .Y(n105) );
  AOI21X4 U334 ( .A0(n149), .A1(n136), .B0(n137), .Y(n135) );
  OAI21X1 U335 ( .A0(n138), .A1(n144), .B0(n139), .Y(n137) );
  NAND2XL U336 ( .A(n212), .B(n154), .Y(n22) );
  NOR2X2 U337 ( .A(n357), .B(n138), .Y(n136) );
  XNOR2X2 U338 ( .A(n92), .B(n11), .Y(SUM[21]) );
  XNOR2X1 U339 ( .A(n38), .B(n2), .Y(SUM[30]) );
  AOI21X1 U340 ( .A0(n38), .A1(n34), .B0(n35), .Y(n33) );
  NAND2X4 U341 ( .A(n367), .B(n40), .Y(n38) );
  NOR2X2 U342 ( .A(n337), .B(A[5]), .Y(n180) );
  BUFX4 U343 ( .A(B[25]), .Y(n330) );
  INVXL U344 ( .A(n118), .Y(n116) );
  INVXL U345 ( .A(n75), .Y(n199) );
  NOR2X4 U346 ( .A(n80), .B(n75), .Y(n73) );
  NOR2X2 U347 ( .A(B[23]), .B(A[23]), .Y(n75) );
  NOR2X2 U348 ( .A(n68), .B(n63), .Y(n61) );
  NOR2X2 U349 ( .A(n321), .B(A[24]), .Y(n68) );
  NOR2X2 U350 ( .A(n330), .B(A[25]), .Y(n63) );
  BUFX3 U351 ( .A(B[4]), .Y(n335) );
  BUFX3 U352 ( .A(B[12]), .Y(n336) );
  BUFX3 U353 ( .A(B[5]), .Y(n337) );
  BUFX4 U354 ( .A(B[7]), .Y(n338) );
  NAND2X1 U355 ( .A(n339), .B(n340), .Y(n341) );
  NAND2X2 U356 ( .A(n341), .B(n151), .Y(n149) );
  NAND2XL U357 ( .A(n322), .B(A[11]), .Y(n151) );
  INVX1 U358 ( .A(n156), .Y(n155) );
  INVXL U359 ( .A(n148), .Y(n146) );
  XNOR2X4 U360 ( .A(n145), .B(n20), .Y(SUM[12]) );
  NAND2X6 U361 ( .A(n369), .B(n72), .Y(n70) );
  NAND2X2 U362 ( .A(n327), .B(n368), .Y(n369) );
  INVXL U363 ( .A(n135), .Y(n346) );
  OR2X8 U364 ( .A(n345), .B(n346), .Y(n133) );
  NAND2X2 U365 ( .A(n148), .B(n136), .Y(n134) );
  INVX3 U366 ( .A(n133), .Y(n132) );
  NAND2X4 U368 ( .A(n362), .B(n48), .Y(n46) );
  AO21X4 U369 ( .A0(n105), .A1(n101), .B0(n102), .Y(n365) );
  AND2X4 U370 ( .A(n156), .B(n107), .Y(n355) );
  NOR2X1 U371 ( .A(n134), .B(n109), .Y(n107) );
  INVXL U372 ( .A(n177), .Y(n176) );
  CLKINVX1 U373 ( .A(n8), .Y(n351) );
  INVXL U374 ( .A(n70), .Y(n350) );
  NAND2XL U375 ( .A(n70), .B(n8), .Y(n352) );
  NAND2X1 U376 ( .A(n321), .B(A[24]), .Y(n69) );
  NAND2X2 U377 ( .A(n336), .B(A[12]), .Y(n144) );
  NOR2X1 U378 ( .A(n336), .B(A[12]), .Y(n143) );
  NAND2X1 U379 ( .A(n338), .B(A[7]), .Y(n170) );
  AND2XL U380 ( .A(n124), .B(n111), .Y(n348) );
  NOR2X4 U381 ( .A(n338), .B(A[7]), .Y(n169) );
  NAND2X1 U382 ( .A(B[8]), .B(A[8]), .Y(n165) );
  NAND2X2 U383 ( .A(n350), .B(n351), .Y(n353) );
  NAND2X2 U384 ( .A(n352), .B(n353), .Y(SUM[24]) );
  NAND2XL U385 ( .A(n198), .B(n69), .Y(n8) );
  OR2X2 U386 ( .A(n360), .B(n361), .Y(n97) );
  CLKINVX1 U387 ( .A(n99), .Y(n361) );
  AND2X2 U388 ( .A(n97), .B(n88), .Y(n354) );
  NOR2X1 U389 ( .A(B[8]), .B(A[8]), .Y(n164) );
  OAI21X4 U390 ( .A0(n177), .A1(n157), .B0(n158), .Y(n156) );
  NAND2X1 U391 ( .A(B[16]), .B(A[16]), .Y(n119) );
  NAND2X1 U392 ( .A(n326), .B(A[26]), .Y(n55) );
  BUFX4 U393 ( .A(n143), .Y(n357) );
  INVXL U394 ( .A(n86), .Y(n84) );
  XOR2X1 U396 ( .A(n95), .B(n12), .Y(SUM[20]) );
  INVXL U397 ( .A(n93), .Y(n202) );
  OR2X4 U398 ( .A(n106), .B(n47), .Y(n362) );
  NOR2X2 U399 ( .A(B[13]), .B(A[13]), .Y(n138) );
  NOR2X2 U400 ( .A(B[17]), .B(A[17]), .Y(n113) );
  NAND2X1 U401 ( .A(n332), .B(A[20]), .Y(n94) );
  NAND2XL U402 ( .A(B[29]), .B(A[29]), .Y(n40) );
  NAND2X1 U403 ( .A(n73), .B(n61), .Y(n59) );
  NAND2X1 U404 ( .A(n57), .B(n49), .Y(n47) );
  NAND2XL U405 ( .A(n328), .B(n45), .Y(n4) );
  XNOR2XL U406 ( .A(n46), .B(n4), .Y(SUM[28]) );
  NAND2X2 U407 ( .A(B[14]), .B(A[14]), .Y(n131) );
  NAND2X2 U408 ( .A(B[18]), .B(A[18]), .Y(n104) );
  NOR2X1 U409 ( .A(B[18]), .B(A[18]), .Y(n103) );
  NOR2X1 U410 ( .A(n326), .B(A[26]), .Y(n54) );
  NOR2X1 U411 ( .A(B[27]), .B(A[27]), .Y(n51) );
  NOR2X1 U412 ( .A(B[3]), .B(A[3]), .Y(n187) );
  NAND2X1 U413 ( .A(n167), .B(n159), .Y(n157) );
  XOR2X1 U414 ( .A(n185), .B(n28), .Y(SUM[4]) );
  INVXL U415 ( .A(n183), .Y(n218) );
  OAI21XL U416 ( .A0(n185), .A1(n183), .B0(n184), .Y(n182) );
  AOI21X1 U417 ( .A0(n46), .A1(n328), .B0(n43), .Y(n41) );
  CLKINVX1 U418 ( .A(n45), .Y(n43) );
  NAND2BXL U419 ( .AN(n189), .B(n190), .Y(n30) );
  INVX1 U420 ( .A(n30), .Y(SUM[2]) );
  NOR2X2 U421 ( .A(n322), .B(A[11]), .Y(n150) );
  INVXL U422 ( .A(n170), .Y(n359) );
  NOR2X1 U423 ( .A(n104), .B(n98), .Y(n360) );
  NAND2X1 U424 ( .A(A[19]), .B(B[19]), .Y(n99) );
  INVXL U425 ( .A(n149), .Y(n147) );
  INVXL U427 ( .A(n186), .Y(n185) );
  CLKINVX1 U428 ( .A(n71), .Y(n368) );
  XNOR2X1 U430 ( .A(n363), .B(n19), .Y(SUM[13]) );
  XOR2X1 U431 ( .A(n364), .B(n5), .Y(SUM[27]) );
  XNOR2X1 U432 ( .A(n365), .B(n13), .Y(SUM[19]) );
  OAI21X1 U433 ( .A0(n166), .A1(n333), .B0(n165), .Y(n163) );
  XNOR2X1 U434 ( .A(n366), .B(n25), .Y(SUM[7]) );
  AO21XL U435 ( .A0(n323), .A1(n172), .B0(n173), .Y(n366) );
  INVXL U436 ( .A(n37), .Y(n35) );
  NOR2X2 U438 ( .A(n130), .B(n125), .Y(n123) );
  NAND2XL U440 ( .A(B[13]), .B(A[13]), .Y(n139) );
  NAND2XL U441 ( .A(B[9]), .B(A[9]), .Y(n162) );
  NAND2XL U442 ( .A(n331), .B(A[21]), .Y(n91) );
  NAND2XL U443 ( .A(B[17]), .B(A[17]), .Y(n114) );
  NAND2XL U444 ( .A(B[27]), .B(A[27]), .Y(n52) );
  NOR2XL U445 ( .A(B[2]), .B(A[2]), .Y(n189) );
  NOR2X1 U446 ( .A(B[30]), .B(A[30]), .Y(n36) );
  INVXL U447 ( .A(n73), .Y(n71) );
  INVX1 U448 ( .A(n74), .Y(n72) );
  AOI21X1 U449 ( .A0(n323), .A1(n167), .B0(n168), .Y(n166) );
  NAND2X1 U450 ( .A(n96), .B(n88), .Y(n86) );
  OAI21XL U451 ( .A0(n63), .A1(n69), .B0(n64), .Y(n62) );
  AOI21X1 U452 ( .A0(n58), .A1(n49), .B0(n50), .Y(n48) );
  NOR2X1 U453 ( .A(n54), .B(n51), .Y(n49) );
  XNOR2X1 U454 ( .A(n323), .B(n26), .Y(SUM[6]) );
  NAND2X1 U455 ( .A(n172), .B(n175), .Y(n26) );
  NAND2X1 U456 ( .A(n195), .B(n52), .Y(n5) );
  OAI21XL U457 ( .A0(n51), .A1(n55), .B0(n52), .Y(n50) );
  XNOR2X1 U458 ( .A(n182), .B(n27), .Y(SUM[5]) );
  NAND2X1 U459 ( .A(n217), .B(n181), .Y(n27) );
  XNOR2X1 U460 ( .A(n163), .B(n23), .Y(SUM[9]) );
  NAND2X1 U461 ( .A(n213), .B(n162), .Y(n23) );
  XNOR2X1 U462 ( .A(n152), .B(n21), .Y(SUM[11]) );
  NAND2X1 U463 ( .A(n339), .B(n151), .Y(n21) );
  NAND2X1 U464 ( .A(n201), .B(n91), .Y(n11) );
  XOR2X1 U465 ( .A(n41), .B(n3), .Y(SUM[29]) );
  NAND2X1 U466 ( .A(n1), .B(n40), .Y(n3) );
  XNOR2X1 U467 ( .A(n120), .B(n16), .Y(SUM[16]) );
  NAND2X1 U468 ( .A(n116), .B(n119), .Y(n16) );
  NAND2X1 U470 ( .A(n205), .B(n114), .Y(n15) );
  NAND2X1 U472 ( .A(n101), .B(n104), .Y(n14) );
  NAND2X1 U473 ( .A(n203), .B(n99), .Y(n13) );
  NAND2X1 U474 ( .A(n202), .B(n94), .Y(n12) );
  XNOR2X1 U475 ( .A(n327), .B(n10), .Y(SUM[22]) );
  NAND2X1 U476 ( .A(n78), .B(n81), .Y(n10) );
  XOR2X1 U477 ( .A(n77), .B(n9), .Y(SUM[23]) );
  NAND2X1 U478 ( .A(n199), .B(n76), .Y(n9) );
  AOI21X1 U479 ( .A0(n327), .A1(n78), .B0(n79), .Y(n77) );
  CLKINVX1 U480 ( .A(n68), .Y(n198) );
  XOR2X1 U481 ( .A(n166), .B(n24), .Y(SUM[8]) );
  NAND2X1 U482 ( .A(n214), .B(n165), .Y(n24) );
  CLKINVX1 U483 ( .A(n333), .Y(n214) );
  XOR2X1 U484 ( .A(n324), .B(n22), .Y(SUM[10]) );
  NAND2X1 U485 ( .A(n141), .B(n144), .Y(n20) );
  XOR2X1 U486 ( .A(n132), .B(n18), .Y(SUM[14]) );
  NAND2X1 U487 ( .A(n128), .B(n131), .Y(n18) );
  NAND2BX1 U488 ( .AN(n36), .B(n37), .Y(n2) );
  CLKINVX1 U489 ( .A(n174), .Y(n172) );
  CLKINVX1 U490 ( .A(n357), .Y(n141) );
  CLKINVX1 U491 ( .A(n130), .Y(n128) );
  CLKINVX1 U492 ( .A(n80), .Y(n78) );
  CLKINVX1 U493 ( .A(n36), .Y(n34) );
  CLKINVX1 U494 ( .A(n69), .Y(n67) );
  NAND2X1 U495 ( .A(n215), .B(n170), .Y(n25) );
  NAND2X1 U496 ( .A(n218), .B(n184), .Y(n28) );
  NAND2X1 U497 ( .A(n209), .B(n139), .Y(n19) );
  XOR2X1 U498 ( .A(n127), .B(n17), .Y(SUM[15]) );
  NAND2X1 U500 ( .A(n197), .B(n64), .Y(n7) );
  CLKINVX1 U501 ( .A(n63), .Y(n197) );
  NAND2X1 U502 ( .A(n196), .B(n55), .Y(n6) );
  CLKINVX1 U503 ( .A(n54), .Y(n196) );
  XOR2X1 U504 ( .A(n29), .B(n190), .Y(SUM[3]) );
  NAND2X1 U505 ( .A(n219), .B(n188), .Y(n29) );
  CLKINVX1 U506 ( .A(n187), .Y(n219) );
  CLKINVX1 U507 ( .A(n175), .Y(n173) );
  CLKINVX1 U508 ( .A(n144), .Y(n142) );
  CLKINVX1 U509 ( .A(n131), .Y(n129) );
  CLKINVX1 U510 ( .A(n119), .Y(n117) );
  CLKINVX1 U511 ( .A(n104), .Y(n102) );
  CLKINVX1 U512 ( .A(n81), .Y(n79) );
  CLKINVX1 U513 ( .A(n51), .Y(n195) );
  CLKINVX1 U514 ( .A(n121), .Y(n217) );
  CLKINVX1 U515 ( .A(n169), .Y(n215) );
  CLKINVX1 U516 ( .A(n161), .Y(n213) );
  CLKINVX1 U517 ( .A(n138), .Y(n209) );
  CLKINVX1 U518 ( .A(n125), .Y(n207) );
  CLKINVX1 U519 ( .A(n113), .Y(n205) );
  CLKINVX1 U520 ( .A(n82), .Y(n203) );
  CLKINVX1 U521 ( .A(n90), .Y(n201) );
  OR2X1 U522 ( .A(B[31]), .B(A[31]), .Y(n370) );
  NAND2X1 U523 ( .A(B[30]), .B(A[30]), .Y(n37) );
  NAND2X1 U524 ( .A(B[28]), .B(A[28]), .Y(n45) );
  NAND2X1 U525 ( .A(B[3]), .B(A[3]), .Y(n188) );
  NAND2X1 U528 ( .A(B[31]), .B(A[31]), .Y(n32) );
  CLKBUFX3 U529 ( .A(A[1]), .Y(SUM[1]) );
  CLKBUFX3 U530 ( .A(A[0]), .Y(SUM[0]) );
  INVXL U1 ( .A(n65), .Y(n1) );
  OAI2BB1X4 U2 ( .A0N(n31), .A1N(n202), .B0(n94), .Y(n92) );
  CLKINVX20 U3 ( .A(n95), .Y(n31) );
  OA21X4 U4 ( .A0(n324), .A1(n153), .B0(n154), .Y(n39) );
  CLKINVX20 U5 ( .A(n39), .Y(n152) );
  OAI2BB1X4 U6 ( .A0N(n105), .A1N(n84), .B0(n87), .Y(n327) );
  XNOR2X4 U7 ( .A(n42), .B(n15), .Y(SUM[17]) );
  AO21X4 U8 ( .A0(n120), .A1(n116), .B0(n117), .Y(n42) );
  NOR2BX4 U9 ( .AN(n44), .B(n97), .Y(n95) );
  NAND2X8 U10 ( .A(n105), .B(n96), .Y(n44) );
  AO21X4 U11 ( .A0(n105), .A1(n57), .B0(n58), .Y(n53) );
  CLKINVX20 U12 ( .A(n53), .Y(n56) );
  OR2X8 U13 ( .A(n66), .B(n65), .Y(n367) );
  CLKINVX20 U14 ( .A(n329), .Y(n65) );
  AOI21X4 U15 ( .A0(n46), .A1(n328), .B0(n43), .Y(n66) );
  CLKBUFX20 U16 ( .A(n98), .Y(n82) );
  XNOR2X4 U17 ( .A(n33), .B(n83), .Y(SUM[31]) );
  CLKAND2X12 U18 ( .A(n370), .B(n32), .Y(n83) );
  XNOR2X4 U19 ( .A(n85), .B(n7), .Y(SUM[25]) );
  AO21X4 U20 ( .A0(n70), .A1(n198), .B0(n67), .Y(n85) );
  NOR2BX4 U21 ( .AN(n337), .B(n115), .Y(n100) );
  CLKINVX20 U22 ( .A(n100), .Y(n181) );
  CLKINVX20 U23 ( .A(A[5]), .Y(n115) );
  CLKBUFX20 U24 ( .A(n180), .Y(n121) );
endmodule


module InstructionDecode_test_1 ( clk, rst, stall, PCadd4, Instruction, 
        PCbranched, Reg_W, WriteData, WB, MEM, EX, RData1, RData2, next_RData1, 
        Immediate_SE, RegisterRd, RegisterRs, RegisterRt, MEM_RegWrite, RegDst, 
        Jump, Branch, MemRead, MemtoReg, MemWrite, ALUOp, ALUSrc, RegWrite, 
        Bubble, PCBuffer_valid, equal, EX_RegWriteData, MEM_RegWriteData, 
        BrForwardA, BrForwardB, PredictMiss, BranchTaken, test_si2, test_si1, 
        test_so2, test_so1, test_se );
  input [31:0] PCadd4;
  input [31:0] Instruction;
  output [31:0] PCbranched;
  input [4:0] Reg_W;
  input [31:0] WriteData;
  output [1:0] WB;
  output [2:0] MEM;
  output [6:0] EX;
  output [31:0] RData1;
  output [31:0] RData2;
  output [31:0] next_RData1;
  output [31:0] Immediate_SE;
  output [4:0] RegisterRd;
  output [4:0] RegisterRs;
  output [4:0] RegisterRt;
  input [2:0] ALUOp;
  input [31:0] EX_RegWriteData;
  input [31:0] MEM_RegWriteData;
  input [1:0] BrForwardA;
  input [1:0] BrForwardB;
  input clk, rst, stall, MEM_RegWrite, RegDst, Jump, Branch, MemRead, MemtoReg,
         MemWrite, ALUSrc, RegWrite, Bubble, BranchTaken, test_si2, test_si1,
         test_se;
  output PCBuffer_valid, equal, PredictMiss, test_so2, test_so1;
  wire   n1941, n1943, n1945, n1947, n1949, n1951, n1953, n1955, n1957, n1959,
         n1961, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26,
         \regfile[15][31] , \regfile[15][30] , \regfile[15][29] ,
         \regfile[15][28] , \regfile[15][27] , \regfile[15][26] ,
         \regfile[15][25] , \regfile[15][24] , \regfile[15][23] ,
         \regfile[15][22] , \regfile[15][21] , \regfile[15][20] ,
         \regfile[15][19] , \regfile[15][18] , \regfile[15][17] ,
         \regfile[15][16] , \regfile[15][15] , \regfile[15][14] ,
         \regfile[15][13] , \regfile[15][12] , \regfile[15][11] ,
         \regfile[15][10] , \regfile[15][9] , \regfile[15][8] ,
         \regfile[15][7] , \regfile[15][6] , \regfile[15][5] ,
         \regfile[15][4] , \regfile[15][3] , \regfile[15][2] ,
         \regfile[15][1] , \regfile[15][0] , \regfile[14][31] ,
         \regfile[14][30] , \regfile[14][29] , \regfile[14][28] ,
         \regfile[14][27] , \regfile[14][26] , \regfile[14][25] ,
         \regfile[14][24] , \regfile[14][23] , \regfile[14][22] ,
         \regfile[14][21] , \regfile[14][20] , \regfile[14][19] ,
         \regfile[14][18] , \regfile[14][17] , \regfile[14][16] ,
         \regfile[14][15] , \regfile[14][14] , \regfile[14][13] ,
         \regfile[14][12] , \regfile[14][11] , \regfile[14][10] ,
         \regfile[14][9] , \regfile[14][8] , \regfile[14][7] ,
         \regfile[14][6] , \regfile[14][5] , \regfile[14][4] ,
         \regfile[14][3] , \regfile[14][2] , \regfile[14][1] ,
         \regfile[14][0] , \regfile[13][31] , \regfile[13][30] ,
         \regfile[13][29] , \regfile[13][28] , \regfile[13][27] ,
         \regfile[13][26] , \regfile[13][25] , \regfile[13][24] ,
         \regfile[13][23] , \regfile[13][22] , \regfile[13][21] ,
         \regfile[13][20] , \regfile[13][19] , \regfile[13][18] ,
         \regfile[13][17] , \regfile[13][16] , \regfile[13][15] ,
         \regfile[13][14] , \regfile[13][13] , \regfile[13][12] ,
         \regfile[13][11] , \regfile[13][10] , \regfile[13][9] ,
         \regfile[13][8] , \regfile[13][7] , \regfile[13][6] ,
         \regfile[13][5] , \regfile[13][4] , \regfile[13][3] ,
         \regfile[13][2] , \regfile[13][1] , \regfile[13][0] ,
         \regfile[12][31] , \regfile[12][30] , \regfile[12][29] ,
         \regfile[12][28] , \regfile[12][27] , \regfile[12][26] ,
         \regfile[12][25] , \regfile[12][24] , \regfile[12][23] ,
         \regfile[12][22] , \regfile[12][21] , \regfile[12][20] ,
         \regfile[12][19] , \regfile[12][18] , \regfile[12][17] ,
         \regfile[12][16] , \regfile[12][15] , \regfile[12][14] ,
         \regfile[12][13] , \regfile[12][12] , \regfile[12][11] ,
         \regfile[12][10] , \regfile[12][9] , \regfile[12][8] ,
         \regfile[12][7] , \regfile[12][6] , \regfile[12][5] ,
         \regfile[12][4] , \regfile[12][3] , \regfile[12][2] ,
         \regfile[12][1] , \regfile[12][0] , \regfile[11][31] ,
         \regfile[11][30] , \regfile[11][29] , \regfile[11][28] ,
         \regfile[11][27] , \regfile[11][26] , \regfile[11][25] ,
         \regfile[11][24] , \regfile[11][23] , \regfile[11][22] ,
         \regfile[11][21] , \regfile[11][20] , \regfile[11][19] ,
         \regfile[11][18] , \regfile[11][17] , \regfile[11][16] ,
         \regfile[11][15] , \regfile[11][14] , \regfile[11][13] ,
         \regfile[11][12] , \regfile[11][11] , \regfile[11][10] ,
         \regfile[11][9] , \regfile[11][8] , \regfile[11][7] ,
         \regfile[11][6] , \regfile[11][5] , \regfile[11][4] ,
         \regfile[11][3] , \regfile[11][2] , \regfile[11][1] ,
         \regfile[11][0] , \regfile[10][31] , \regfile[10][30] ,
         \regfile[10][29] , \regfile[10][28] , \regfile[10][27] ,
         \regfile[10][26] , \regfile[10][25] , \regfile[10][24] ,
         \regfile[10][23] , \regfile[10][22] , \regfile[10][21] ,
         \regfile[10][20] , \regfile[10][19] , \regfile[10][18] ,
         \regfile[10][17] , \regfile[10][16] , \regfile[10][15] ,
         \regfile[10][14] , \regfile[10][13] , \regfile[10][12] ,
         \regfile[10][11] , \regfile[10][10] , \regfile[10][9] ,
         \regfile[10][8] , \regfile[10][7] , \regfile[10][6] ,
         \regfile[10][5] , \regfile[10][4] , \regfile[10][3] ,
         \regfile[10][2] , \regfile[10][1] , \regfile[10][0] ,
         \regfile[9][31] , \regfile[9][30] , \regfile[9][29] ,
         \regfile[9][28] , \regfile[9][27] , \regfile[9][26] ,
         \regfile[9][25] , \regfile[9][24] , \regfile[9][23] ,
         \regfile[9][22] , \regfile[9][21] , \regfile[9][20] ,
         \regfile[9][19] , \regfile[9][18] , \regfile[9][17] ,
         \regfile[9][16] , \regfile[9][15] , \regfile[9][14] ,
         \regfile[9][13] , \regfile[9][12] , \regfile[9][11] ,
         \regfile[9][10] , \regfile[9][9] , \regfile[9][8] , \regfile[9][7] ,
         \regfile[9][6] , \regfile[9][5] , \regfile[9][4] , \regfile[9][3] ,
         \regfile[9][2] , \regfile[9][1] , \regfile[9][0] , \regfile[8][31] ,
         \regfile[8][30] , \regfile[8][29] , \regfile[8][28] ,
         \regfile[8][27] , \regfile[8][26] , \regfile[8][25] ,
         \regfile[8][24] , \regfile[8][23] , \regfile[8][22] ,
         \regfile[8][21] , \regfile[8][20] , \regfile[8][19] ,
         \regfile[8][18] , \regfile[8][17] , \regfile[8][16] ,
         \regfile[8][15] , \regfile[8][14] , \regfile[8][13] ,
         \regfile[8][12] , \regfile[8][11] , \regfile[8][10] , \regfile[8][9] ,
         \regfile[8][8] , \regfile[8][7] , \regfile[8][6] , \regfile[8][5] ,
         \regfile[8][4] , \regfile[8][3] , \regfile[8][2] , \regfile[8][1] ,
         \regfile[8][0] , \regfile[7][31] , \regfile[7][30] , \regfile[7][29] ,
         \regfile[7][28] , \regfile[7][27] , \regfile[7][26] ,
         \regfile[7][25] , \regfile[7][24] , \regfile[7][23] ,
         \regfile[7][22] , \regfile[7][21] , \regfile[7][20] ,
         \regfile[7][19] , \regfile[7][18] , \regfile[7][17] ,
         \regfile[7][16] , \regfile[7][15] , \regfile[7][14] ,
         \regfile[7][13] , \regfile[7][12] , \regfile[7][11] ,
         \regfile[7][10] , \regfile[7][9] , \regfile[7][8] , \regfile[7][7] ,
         \regfile[7][6] , \regfile[7][5] , \regfile[7][4] , \regfile[7][3] ,
         \regfile[7][2] , \regfile[7][1] , \regfile[7][0] , \regfile[6][31] ,
         \regfile[6][30] , \regfile[6][29] , \regfile[6][28] ,
         \regfile[6][27] , \regfile[6][26] , \regfile[6][25] ,
         \regfile[6][24] , \regfile[6][23] , \regfile[6][22] ,
         \regfile[6][21] , \regfile[6][20] , \regfile[6][19] ,
         \regfile[6][18] , \regfile[6][17] , \regfile[6][16] ,
         \regfile[6][15] , \regfile[6][14] , \regfile[6][13] ,
         \regfile[6][12] , \regfile[6][11] , \regfile[6][10] , \regfile[6][9] ,
         \regfile[6][8] , \regfile[6][7] , \regfile[6][6] , \regfile[6][5] ,
         \regfile[6][4] , \regfile[6][3] , \regfile[6][2] , \regfile[6][1] ,
         \regfile[6][0] , \regfile[5][31] , \regfile[5][30] , \regfile[5][29] ,
         \regfile[5][28] , \regfile[5][27] , \regfile[5][26] ,
         \regfile[5][25] , \regfile[5][24] , \regfile[5][23] ,
         \regfile[5][22] , \regfile[5][21] , \regfile[5][20] ,
         \regfile[5][19] , \regfile[5][18] , \regfile[5][17] ,
         \regfile[5][16] , \regfile[5][15] , \regfile[5][14] ,
         \regfile[5][13] , \regfile[5][12] , \regfile[5][11] ,
         \regfile[5][10] , \regfile[5][9] , \regfile[5][8] , \regfile[5][7] ,
         \regfile[5][6] , \regfile[5][5] , \regfile[5][4] , \regfile[5][3] ,
         \regfile[5][2] , \regfile[5][1] , \regfile[5][0] , \regfile[4][31] ,
         \regfile[4][30] , \regfile[4][29] , \regfile[4][28] ,
         \regfile[4][27] , \regfile[4][26] , \regfile[4][25] ,
         \regfile[4][24] , \regfile[4][23] , \regfile[4][22] ,
         \regfile[4][21] , \regfile[4][20] , \regfile[4][19] ,
         \regfile[4][18] , \regfile[4][17] , \regfile[4][16] ,
         \regfile[4][15] , \regfile[4][14] , \regfile[4][13] ,
         \regfile[4][12] , \regfile[4][11] , \regfile[4][10] , \regfile[4][9] ,
         \regfile[4][8] , \regfile[4][7] , \regfile[4][6] , \regfile[4][5] ,
         \regfile[4][4] , \regfile[4][3] , \regfile[4][2] , \regfile[4][1] ,
         \regfile[4][0] , \regfile[3][31] , \regfile[3][30] , \regfile[3][29] ,
         \regfile[3][28] , \regfile[3][27] , \regfile[3][26] ,
         \regfile[3][25] , \regfile[3][24] , \regfile[3][22] ,
         \regfile[3][21] , \regfile[3][17] , \regfile[3][16] ,
         \regfile[3][15] , \regfile[3][14] , \regfile[3][13] ,
         \regfile[3][12] , \regfile[3][11] , \regfile[3][9] , \regfile[3][8] ,
         \regfile[3][6] , \regfile[3][5] , \regfile[3][3] , \regfile[3][2] ,
         \regfile[3][1] , \regfile[1][31] , \regfile[1][30] , \regfile[1][29] ,
         \regfile[1][28] , \regfile[1][27] , \regfile[1][26] ,
         \regfile[1][25] , \regfile[1][24] , \regfile[1][23] ,
         \regfile[1][22] , \regfile[1][21] , \regfile[1][20] ,
         \regfile[1][19] , \regfile[1][18] , \regfile[1][17] ,
         \regfile[1][16] , \regfile[1][15] , \regfile[1][14] ,
         \regfile[1][13] , \regfile[1][12] , \regfile[1][11] ,
         \regfile[1][10] , \regfile[1][9] , \regfile[1][8] , \regfile[1][7] ,
         \regfile[1][6] , \regfile[1][5] , \regfile[1][4] , \regfile[1][3] ,
         \regfile[1][2] , \regfile[1][1] , \regfile[1][0] , \regfile[31][31] ,
         \regfile[31][30] , \regfile[31][29] , \regfile[31][28] ,
         \regfile[31][27] , \regfile[31][26] , \regfile[31][25] ,
         \regfile[31][24] , \regfile[31][23] , \regfile[31][22] ,
         \regfile[31][21] , \regfile[31][20] , \regfile[31][19] ,
         \regfile[31][18] , \regfile[31][17] , \regfile[31][16] ,
         \regfile[31][15] , \regfile[31][14] , \regfile[31][13] ,
         \regfile[31][12] , \regfile[31][11] , \regfile[31][10] ,
         \regfile[31][9] , \regfile[31][8] , \regfile[31][7] ,
         \regfile[31][6] , \regfile[31][5] , \regfile[31][4] ,
         \regfile[31][3] , \regfile[31][2] , \regfile[31][1] ,
         \regfile[31][0] , \regfile[30][31] , \regfile[30][30] ,
         \regfile[30][29] , \regfile[30][28] , \regfile[30][27] ,
         \regfile[30][26] , \regfile[30][25] , \regfile[30][24] ,
         \regfile[30][23] , \regfile[30][22] , \regfile[30][21] ,
         \regfile[30][20] , \regfile[30][19] , \regfile[30][18] ,
         \regfile[30][17] , \regfile[30][16] , \regfile[30][15] ,
         \regfile[30][14] , \regfile[30][13] , \regfile[30][12] ,
         \regfile[30][11] , \regfile[30][10] , \regfile[30][9] ,
         \regfile[30][8] , \regfile[30][7] , \regfile[30][6] ,
         \regfile[30][5] , \regfile[30][4] , \regfile[30][3] ,
         \regfile[30][2] , \regfile[30][1] , \regfile[30][0] ,
         \regfile[29][31] , \regfile[29][30] , \regfile[29][29] ,
         \regfile[29][28] , \regfile[29][27] , \regfile[29][26] ,
         \regfile[29][25] , \regfile[29][24] , \regfile[29][23] ,
         \regfile[29][22] , \regfile[29][21] , \regfile[29][20] ,
         \regfile[29][19] , \regfile[29][18] , \regfile[29][17] ,
         \regfile[29][16] , \regfile[29][15] , \regfile[29][14] ,
         \regfile[29][13] , \regfile[29][12] , \regfile[29][11] ,
         \regfile[29][10] , \regfile[29][9] , \regfile[29][8] ,
         \regfile[29][7] , \regfile[29][6] , \regfile[29][5] ,
         \regfile[29][4] , \regfile[29][3] , \regfile[29][2] ,
         \regfile[29][1] , \regfile[29][0] , \regfile[28][31] ,
         \regfile[28][30] , \regfile[28][29] , \regfile[28][28] ,
         \regfile[28][27] , \regfile[28][26] , \regfile[28][25] ,
         \regfile[28][24] , \regfile[28][23] , \regfile[28][22] ,
         \regfile[28][21] , \regfile[28][20] , \regfile[28][19] ,
         \regfile[28][18] , \regfile[28][17] , \regfile[28][16] ,
         \regfile[28][15] , \regfile[28][14] , \regfile[28][13] ,
         \regfile[28][12] , \regfile[28][11] , \regfile[28][10] ,
         \regfile[28][9] , \regfile[28][8] , \regfile[28][7] ,
         \regfile[28][6] , \regfile[28][5] , \regfile[28][4] ,
         \regfile[28][3] , \regfile[28][2] , \regfile[28][1] ,
         \regfile[28][0] , \regfile[27][31] , \regfile[27][30] ,
         \regfile[27][29] , \regfile[27][28] , \regfile[27][27] ,
         \regfile[27][26] , \regfile[27][25] , \regfile[27][24] ,
         \regfile[27][23] , \regfile[27][22] , \regfile[27][21] ,
         \regfile[27][20] , \regfile[27][19] , \regfile[27][18] ,
         \regfile[27][17] , \regfile[27][16] , \regfile[27][15] ,
         \regfile[27][14] , \regfile[27][13] , \regfile[27][12] ,
         \regfile[27][11] , \regfile[27][10] , \regfile[27][9] ,
         \regfile[27][8] , \regfile[27][7] , \regfile[27][6] ,
         \regfile[27][5] , \regfile[27][4] , \regfile[27][3] ,
         \regfile[27][2] , \regfile[27][1] , \regfile[27][0] ,
         \regfile[26][31] , \regfile[26][30] , \regfile[26][29] ,
         \regfile[26][28] , \regfile[26][27] , \regfile[26][26] ,
         \regfile[26][25] , \regfile[26][24] , \regfile[26][23] ,
         \regfile[26][22] , \regfile[26][21] , \regfile[26][20] ,
         \regfile[26][19] , \regfile[26][18] , \regfile[26][17] ,
         \regfile[26][16] , \regfile[26][15] , \regfile[26][14] ,
         \regfile[26][13] , \regfile[26][12] , \regfile[26][11] ,
         \regfile[26][10] , \regfile[26][9] , \regfile[26][8] ,
         \regfile[26][7] , \regfile[26][6] , \regfile[26][5] ,
         \regfile[26][4] , \regfile[26][3] , \regfile[26][2] ,
         \regfile[26][1] , \regfile[26][0] , \regfile[25][31] ,
         \regfile[25][30] , \regfile[25][29] , \regfile[25][28] ,
         \regfile[25][27] , \regfile[25][26] , \regfile[25][25] ,
         \regfile[25][24] , \regfile[25][23] , \regfile[25][22] ,
         \regfile[25][21] , \regfile[25][20] , \regfile[25][19] ,
         \regfile[25][18] , \regfile[25][17] , \regfile[25][16] ,
         \regfile[25][15] , \regfile[25][14] , \regfile[25][13] ,
         \regfile[25][12] , \regfile[25][11] , \regfile[25][10] ,
         \regfile[25][9] , \regfile[25][8] , \regfile[25][7] ,
         \regfile[25][6] , \regfile[25][5] , \regfile[25][4] ,
         \regfile[25][3] , \regfile[25][2] , \regfile[25][1] ,
         \regfile[25][0] , \regfile[24][31] , \regfile[24][30] ,
         \regfile[24][29] , \regfile[24][28] , \regfile[24][27] ,
         \regfile[24][26] , \regfile[24][25] , \regfile[24][24] ,
         \regfile[24][23] , \regfile[24][22] , \regfile[24][21] ,
         \regfile[24][20] , \regfile[24][19] , \regfile[24][18] ,
         \regfile[24][17] , \regfile[24][16] , \regfile[24][15] ,
         \regfile[24][14] , \regfile[24][13] , \regfile[24][12] ,
         \regfile[24][11] , \regfile[24][10] , \regfile[24][9] ,
         \regfile[24][8] , \regfile[24][7] , \regfile[24][6] ,
         \regfile[24][5] , \regfile[24][4] , \regfile[24][3] ,
         \regfile[24][2] , \regfile[24][1] , \regfile[24][0] ,
         \regfile[23][31] , \regfile[23][30] , \regfile[23][29] ,
         \regfile[23][28] , \regfile[23][27] , \regfile[23][26] ,
         \regfile[23][25] , \regfile[23][24] , \regfile[23][23] ,
         \regfile[23][22] , \regfile[23][21] , \regfile[23][20] ,
         \regfile[23][19] , \regfile[23][18] , \regfile[23][17] ,
         \regfile[23][16] , \regfile[23][15] , \regfile[23][14] ,
         \regfile[23][13] , \regfile[23][12] , \regfile[23][11] ,
         \regfile[23][10] , \regfile[23][9] , \regfile[23][8] ,
         \regfile[23][7] , \regfile[23][6] , \regfile[23][5] ,
         \regfile[23][4] , \regfile[23][3] , \regfile[23][2] ,
         \regfile[23][1] , \regfile[23][0] , \regfile[22][31] ,
         \regfile[22][30] , \regfile[22][29] , \regfile[22][28] ,
         \regfile[22][27] , \regfile[22][26] , \regfile[22][25] ,
         \regfile[22][24] , \regfile[22][23] , \regfile[22][22] ,
         \regfile[22][21] , \regfile[22][20] , \regfile[22][19] ,
         \regfile[22][18] , \regfile[22][17] , \regfile[22][16] ,
         \regfile[22][15] , \regfile[22][14] , \regfile[22][13] ,
         \regfile[22][12] , \regfile[22][11] , \regfile[22][10] ,
         \regfile[22][9] , \regfile[22][8] , \regfile[22][7] ,
         \regfile[22][6] , \regfile[22][5] , \regfile[22][4] ,
         \regfile[22][3] , \regfile[22][2] , \regfile[22][1] ,
         \regfile[22][0] , \regfile[21][31] , \regfile[21][30] ,
         \regfile[21][29] , \regfile[21][28] , \regfile[21][27] ,
         \regfile[21][26] , \regfile[21][25] , \regfile[21][24] ,
         \regfile[21][23] , \regfile[21][22] , \regfile[21][21] ,
         \regfile[21][20] , \regfile[21][19] , \regfile[21][18] ,
         \regfile[21][17] , \regfile[21][16] , \regfile[21][15] ,
         \regfile[21][14] , \regfile[21][13] , \regfile[21][12] ,
         \regfile[21][11] , \regfile[21][10] , \regfile[21][9] ,
         \regfile[21][8] , \regfile[21][7] , \regfile[21][6] ,
         \regfile[21][5] , \regfile[21][4] , \regfile[21][3] ,
         \regfile[21][2] , \regfile[21][1] , \regfile[21][0] ,
         \regfile[20][31] , \regfile[20][30] , \regfile[20][29] ,
         \regfile[20][28] , \regfile[20][27] , \regfile[20][26] ,
         \regfile[20][25] , \regfile[20][24] , \regfile[20][23] ,
         \regfile[20][22] , \regfile[20][21] , \regfile[20][20] ,
         \regfile[20][19] , \regfile[20][18] , \regfile[20][17] ,
         \regfile[20][16] , \regfile[20][15] , \regfile[20][14] ,
         \regfile[20][13] , \regfile[20][12] , \regfile[20][11] ,
         \regfile[20][10] , \regfile[20][9] , \regfile[20][8] ,
         \regfile[20][7] , \regfile[20][6] , \regfile[20][5] ,
         \regfile[20][4] , \regfile[20][3] , \regfile[20][2] ,
         \regfile[20][1] , \regfile[20][0] , \regfile[19][31] ,
         \regfile[19][30] , \regfile[19][29] , \regfile[19][28] ,
         \regfile[19][27] , \regfile[19][26] , \regfile[19][25] ,
         \regfile[19][24] , \regfile[19][23] , \regfile[19][22] ,
         \regfile[19][21] , \regfile[19][20] , \regfile[19][19] ,
         \regfile[19][18] , \regfile[19][17] , \regfile[19][16] ,
         \regfile[19][15] , \regfile[19][14] , \regfile[19][13] ,
         \regfile[19][12] , \regfile[19][11] , \regfile[19][10] ,
         \regfile[19][9] , \regfile[19][8] , \regfile[19][7] ,
         \regfile[19][6] , \regfile[19][5] , \regfile[19][4] ,
         \regfile[19][3] , \regfile[19][2] , \regfile[19][1] ,
         \regfile[19][0] , \regfile[18][31] , \regfile[18][30] ,
         \regfile[18][29] , \regfile[18][28] , \regfile[18][27] ,
         \regfile[18][26] , \regfile[18][25] , \regfile[18][24] ,
         \regfile[18][23] , \regfile[18][22] , \regfile[18][21] ,
         \regfile[18][20] , \regfile[18][19] , \regfile[18][18] ,
         \regfile[18][17] , \regfile[18][16] , \regfile[18][15] ,
         \regfile[18][14] , \regfile[18][13] , \regfile[18][12] ,
         \regfile[18][11] , \regfile[18][10] , \regfile[18][9] ,
         \regfile[18][8] , \regfile[18][7] , \regfile[18][6] ,
         \regfile[18][5] , \regfile[18][4] , \regfile[18][3] ,
         \regfile[18][2] , \regfile[18][1] , \regfile[18][0] ,
         \regfile[17][31] , \regfile[17][30] , \regfile[17][29] ,
         \regfile[17][28] , \regfile[17][27] , \regfile[17][26] ,
         \regfile[17][25] , \regfile[17][24] , \regfile[17][23] ,
         \regfile[17][22] , \regfile[17][21] , \regfile[17][20] ,
         \regfile[17][19] , \regfile[17][18] , \regfile[17][17] ,
         \regfile[17][16] , \regfile[17][15] , \regfile[17][14] ,
         \regfile[17][13] , \regfile[17][12] , \regfile[17][11] ,
         \regfile[17][10] , \regfile[17][9] , \regfile[17][8] ,
         \regfile[17][7] , \regfile[17][6] , \regfile[17][5] ,
         \regfile[17][4] , \regfile[17][3] , \regfile[17][2] ,
         \regfile[17][1] , \regfile[17][0] , \regfile[16][31] ,
         \regfile[16][30] , \regfile[16][29] , \regfile[16][28] ,
         \regfile[16][27] , \regfile[16][26] , \regfile[16][25] ,
         \regfile[16][24] , \regfile[16][23] , \regfile[16][22] ,
         \regfile[16][21] , \regfile[16][20] , \regfile[16][19] ,
         \regfile[16][18] , \regfile[16][17] , \regfile[16][16] ,
         \regfile[16][15] , \regfile[16][14] , \regfile[16][13] ,
         \regfile[16][12] , \regfile[16][11] , \regfile[16][10] ,
         \regfile[16][9] , \regfile[16][8] , \regfile[16][7] ,
         \regfile[16][6] , \regfile[16][5] , \regfile[16][4] ,
         \regfile[16][3] , \regfile[16][2] , \regfile[16][1] ,
         \regfile[16][0] , N116, N117, N118, N119, N120, N121, N122, N123,
         N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134,
         N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145,
         N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156,
         N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, n10, n12, n53, n54, n57, n61, n62, n65, n66, n73, n76, n83, n86,
         n93, n97, n104, n107, n117, n124, n132, n133, n134, n167, n168, n169,
         n170, n172, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n191, n192, n224, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n624, n625, n626, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1614, n1616, n1618, n1620,
         n1622, n1624, n1626, n1628, n1630, n1632, n1634, n1636, n1638, n1640,
         n1642, n1644, n1646, n1648, n1650, n1652, n1654, n1656, n1658, n1660,
         n1662, n1664, n1666, n1668, n1670, n1672, n1674, n1676, n1678, n1680,
         n1682, n1684, n1686, n1688, n1690, n1692, n1694, n1696, n1698, n1700,
         n1702, n1704, n1706, n1708, n1710, n1712, n1714, n1716, n1718, n1720,
         n1722, n1724, n1726, n1728, n1730, n1732, n1734, n1736, n1738, n1740,
         n1742, n1744, n1746, n1748, n1750, n1752, n1754, n1756, n1758, n1760,
         n1762, n1764, n1766, n1768, n1770, n1772, n1774, n1776, n1778, n1780,
         n1782, n1784, n1786, n1788, n1790, n1792, n1794, n1796, n1798, n1800,
         n1802, n1804, n1806, n1808, n1810, n1812, n1814, n1816, n1818, n1820,
         n1822, n1824, n1826, n1828, n1830, n1832, n1834, n1836, n1838, n1840,
         n1842, n1844, n1846, n1848, n1850, n1852, n1854, n1856, n1858, n1860,
         n1862, n1864, n1866, n1868, n1870, n1872, n1874, n1876, n1878, n1880,
         n1882, n1884, n1886, n1888, n1890, n1892, n1894, n1896, n1898, n1900,
         n1902, n1904, n1906, n1908, n1910, n1912, n1914, n1916, n1918, n1920,
         n1922, n1924, n1926, n1928, n1930, n1932, n1934, n1936, n1938, n1940,
         n1942, n1944, n1946, n1948, n1950, n1952, n1954, n1956, n1958, n1960,
         n1962, n1964, n1966, n1968, n1970, n1972, n1974, n1976, n1978, n1980,
         n1982, n1984, n1986, n1988, n1990, n1992, n1994, n1996, n1998, n2000,
         n2002, n2004, n2006, n2008, n2010, n2012, n2014, n2016, n2018, n2020,
         n2022, n2024, n2026, n2028, n2030, n2032, n2034, n2036, n2038, n2040,
         n2042, n2044, n2046, n2048, n2050, n2052, n2054, n2056, n2058, n2060,
         n2062, n2064, n2066, n2068, n2070, n2072, n2074, n2076, n2078, n2080,
         n2082, n2084, n2086, n2088, n2090, n2092, n2094, n2096, n2098, n2100,
         n2102, n2104, n2106, n2108, n2110, n2112, n2114, n2116, n2118, n2120,
         n2122, n2124, n2126, n2128, n2130, n2132, n2134, n2136, n2138, n2140,
         n2142, n2144, n2146, n2148, n2150, n2152, n2154, n2156, n2158, n2160,
         n2162, n2164, n2166, n2168, n2170, n2172, n2174, n2176, n2178, n2180,
         n2182, n2184, n2186, n2188, n2190, n2192, n2194, n2196, n2198, n2200,
         n2202, n2204, n2206, n2208, n2210, n2212, n2214, n2216, n2218, n2220,
         n2222, n2224, n2226, n2228, n2230, n2232, n2234, n2236, n2238, n2240,
         n2242, n2244, n2246, n2248, n2250, n2252, n2254, n2256, n2258, n2260,
         n2262, n2264, n2266, n2268, n2270, n2272, n2274, n2276, n2278, n2280,
         n2282, n2284, n2286, n2288, n2290, n2292, n2294, n2296, n2298, n2300,
         n2302, n2304, n2306, n2308, n2310, n2312, n2314, n2316, n2318, n2320,
         n2322, n2324, n2326, n2328, n2330, n2332, n2334, n2336, n2338, n2340,
         n2342, n2344, n2346, n2348, n2350, n2352, n2354, n2356, n2358, n2360,
         n2362, n2364, n2366, n2368, n2370, n2372, n2374, n2376, n2378, n2380,
         n2382, n2384, n2386, n2388, n2390, n2392, n2394, n2396, n2398, n2400,
         n2402, n2404, n2406, n2408, n2410, n2412, n2414, n2416, n2418, n2420,
         n2422, n2424, n2426, n2428, n2430, n2432, n2434, n2436, n2438, n2440,
         n2442, n2444, n2446, n2448, n2450, n2452, n2454, n2456, n2458, n2460,
         n2462, n2464, n2466, n2468, n2470, n2472, n2474, n2476, n2478, n2480,
         n2482, n2484, n2486, n2488, n2490, n2492, n2494, n2496, n2498, n2500,
         n2502, n2504, n2506, n2508, n2510, n2512, n2514, n2516, n2518, n2520,
         n2522, n2524, n2526, n2528, n2530, n2532, n2534, n2536, n2538, n2540,
         n2542, n2544, n2546, n2548, n2550, n2552, n2554, n2556, n2558, n2560,
         n2562, n2564, n2566, n2568, n2570, n2572, n2574, n2576, n2578, n2580,
         n2582, n2584, n2586, n2588, n2590, n2592, n2594, n2596, n2598, n2600,
         n2602, n2604, n2606, n2608, n2610, n2612, n2614, n2616, n2618, n2620,
         n2622, n2624, n2626, n2628, n2630, n2632, n2634, n2636, n2638, n2640,
         n2642, n2644, n2646, n2648, n2650, n2652, n2654, n2656, n2658, n2660,
         n2662, n2664, n2666, n2668, n2670, n2672, n2674, n2676, n2678, n2680,
         n2682, n2684, n2686, n2688, n2690, n2692, n2694, n2696, n2698, n2700,
         n2702, n2704, n2706, n2708, n2710, n2712, n2714, n2716, n2718, n2720,
         n2722, n2724, n2726, n2728, n2730, n2732, n2734, n2736, n2738, n2740,
         n2742, n2744, n2746, n2748, n2750, n2752, n2754, n2756, n2758, n2760,
         n2762, n2764, n2766, n2768, n2770, n2772, n2774, n2776, n2778, n2780,
         n2782, n2784, n2786, n2788, n2790, n2792, n2794, n2796, n2798, n2800,
         n2802, n2804, n2806, n2808, n2810, n2812, n2814, n2816, n2818, n2820,
         n2822, n2824, n2826, n2828, n2830, n2832, n2834, n2836, n2838, n2840,
         n2842, n2844, n2846, n2848, n2850, n2852, n2854, n2856, n2858, n2860,
         n2862, n2864, n2866, n2868, n2870, n2872, n2874, n2876, n2878, n2880,
         n2882, n2884, n2886, n2888, n2890, n2892, n2894, n2896, n2898, n2900,
         n2902, n2904, n2906, n2908, n2910, n2912, n2914, n2916, n2918, n2920,
         n2922, n2924, n2926, n2928, n2930, n2932, n2934, n2936, n2938, n2940,
         n2942, n2944, n2946, n2948, n2950, n2952, n2954, n2956, n2958, n2960,
         n2962, n2964, n2966, n2968, n2970, n2972, n2974, n2976, n2978, n2980,
         n2982, n2984, n2986, n2988, n2990, n2992, n2994, n2996, n2998, n3000,
         n3002, n3004, n3006, n3008, n3010, n3012, n3014, n3016, n3018, n3020,
         n3022, n3024, n3026, n3028, n3030, n3032, n3034, n3036, n3038, n3040,
         n3042, n3044, n3046, n3048, n3050, n3052, n3054, n3056, n3058, n3060,
         n3062, n3064, n3066, n3068, n3070, n3072, n3074, n3076, n3078, n3080,
         n3082, n3084, n3086, n3088, n3090, n3092, n3094, n3096, n3098, n3100,
         n3102, n3104, n3106, n3108, n3110, n3112, n3114, n3116, n3118, n3120,
         n3122, n3124, n3126, n3128, n3130, n3132, n3134, n3136, n3138, n3140,
         n3142, n3144, n3146, n3148, n3150, n3152, n3154, n3156, n3158, n3160,
         n3162, n3164, n3166, n3168, n3170, n3172, n3174, n3176, n3178, n3180,
         n3182, n3184, n3186, n3188, n3190, n3192, n3194, n3196, n3198, n3200,
         n3202, n3204, n3206, n3208, n3210, n3212, n3214, n3216, n3218, n3220,
         n3222, n3224, n3226, n3228, n3230, n3232, n3234, n3236, n3238, n3240,
         n3242, n3244, n3246, n3248, n3250, n3252, n3254, n3256, n3258, n3260,
         n3262, n3264, n3266, n3268, n3270, n3272, n3274, n3276, n3278, n3280,
         n3282, n3284, n3286, n3288, n3290, n3292, n3294, n3296, n3298, n3300,
         n3302, n3304, n3306, n3308, n3310, n3312, n3314, n3316, n3318, n3320,
         n3322, n3324, n3326, n3328, n3330, n3332, n3334, n3336, n3338, n3340,
         n3342, n3344, n3346, n3348, n3350, n3352, n3354, n3356, n3358, n3360,
         n3362, n3364, n3366, n3368, n3370, n3372, n3374, n3376, n3378, n3380,
         n3382, n3384, n3386, n3388, n3390, n3392, n3394, n3396, n3398, n3400,
         n3402, n3404, n3406, n3408, n3410, n3412, n3414, n3416, n3418, n3420,
         n3422, n3424, n3426, n3428, n3430, n3432, n3434, n3436, n3438, n3440,
         n3442, n3444, n3446, n3448, n3450, n3452, n3454, n3456, n3458, n3460,
         n3462, n3464, n3466, n3468, n3470, n3472, n3474, n3476, n3478, n3480,
         n3482, n3484, n3486, n3488, n3490, n3492, n3494, n3496, n3498, n3500,
         n3502, n3504, n3506, n3508, n3510, n3512, n3514, n3516, n3518, n3520,
         n3522, n3524, n3526, n3528, n3530, n3532, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, N484, N483, N482, N481, N480, N479, N478, N477, N476,
         N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465,
         N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n11, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n85, n87, n88, n89, n90, n91, n92, n94, n95, n96, n99, n100, n102,
         n103, n105, n106, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n118, n119, n120, n121, n122, n123, n125, n126, n127, n128,
         n129, n130, n131, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n173, n174, n175, n188, n189, n190, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n623, n627, n628,
         n629, n630, n1677, n1679, n1681, n1683, n1685, n1687, n1689, n1691,
         n1693, n1695, n1697, n1699, n1701, n1703, n1705, n1707, n1709, n1711,
         n1713, n1715, n1717, n1719, n1721, n1723, n1725, n1727, n1729, n1731,
         n1733, n1735, n1737, n1739, n1741, n1747, n1749, n1755, n1761, n1777,
         n1779, n1781, n1787, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3799,
         n3800, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4901, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1,
         SYNOPSYS_UNCONNECTED__2, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n55, n56, n58, n59, n60, n63, n64,
         n67, n68, n69, n70, n71, n72, n74, n75, n77, n78, n79, n80, n81, n82,
         n84, n101, n1613, n1615, n1617, n1619, n1621, n1623, n1625, n1627,
         n1629, n1631, n1633, n1635, n1637, n1639, n1641, n1643, n1645, n1647,
         n1649, n1651, n1653, n1655, n1657, n1659, n1661, n1663, n1665, n1667,
         n1669, n1671, n1673, n1675, n1743, n1751, n1753, n1757, n1759, n1763,
         n1765, n1767, n1769, n1771, n1773, n1775, n1783, n1785, n1789, n1791,
         n1793, n1795, n1797, n1799, n1801, n1803, n1805, n1807, n1809, n1811,
         n1813, n1815, n1817, n1819, n1821, n1823, n1825, n1827, n1829, n1831,
         n1833, n1835, n1837, n1839, n1841, n1843, n1845, n1847, n1849, n1851,
         n1853, n1855, n1857, n1859, n1861, n1863, n1865, n1867, n1869, n1871,
         n1873, n1875, n1877, n1879, n1881, n1883, n1885, n1887, n1889, n1891,
         n1893, n1895, n1897, n1899, n1901, n1911, n1913, n1915, n1929, n1931,
         n1935, n1937, n1939;
  wire   [31:0] next_RData2;
  wire   [29:0] next_Immediate_SE;
  assign MEM[2] = 1'b0;
  assign N17 = Instruction[21];
  assign N18 = Instruction[22];
  assign N19 = Instruction[23];
  assign N20 = Instruction[24];
  assign N21 = Instruction[25];
  assign N22 = Instruction[16];
  assign N23 = Instruction[17];
  assign N24 = Instruction[18];
  assign N25 = Instruction[19];
  assign N26 = Instruction[20];
  assign test_so1 = n569;

  XNOR2X2 U5 ( .A(n4848), .B(n4847), .Y(n4849) );
  OAI221X4 U6 ( .A0(n4406), .A1(n4846), .B0(n4841), .B1(n4405), .C0(n4840), 
        .Y(n4848) );
  XNOR2X2 U7 ( .A(n4879), .B(n4878), .Y(n4890) );
  OAI221X4 U8 ( .A0(n4406), .A1(n4877), .B0(n4872), .B1(n4405), .C0(n4871), 
        .Y(n4879) );
  INVX1 U9 ( .A(next_RData1[29]), .Y(n4677) );
  XNOR2X4 U11 ( .A(n4795), .B(n4794), .Y(n4806) );
  OAI221X4 U12 ( .A0(n4416), .A1(n4793), .B0(n4792), .B1(n4413), .C0(n4791), 
        .Y(n4794) );
  INVX4 U14 ( .A(next_RData1[25]), .Y(n4717) );
  OAI221X2 U15 ( .A0(n4407), .A1(n4828), .B0(n4823), .B1(n4405), .C0(n4822), 
        .Y(n4830) );
  INVX1 U16 ( .A(next_RData1[15]), .Y(n4823) );
  OAI221X2 U17 ( .A0(n4406), .A1(n4868), .B0(n4863), .B1(n4405), .C0(n4862), 
        .Y(n4870) );
  OAI221X4 U18 ( .A0(n4407), .A1(n4793), .B0(n4788), .B1(n4405), .C0(n4787), 
        .Y(n4795) );
  XNOR2X2 U19 ( .A(n4957), .B(n4956), .Y(n4976) );
  OAI221X2 U20 ( .A0(n4406), .A1(n4955), .B0(n4950), .B1(n4405), .C0(n4949), 
        .Y(n4957) );
  INVX4 U21 ( .A(next_RData2[0]), .Y(n4954) );
  OAI221X2 U22 ( .A0(n4415), .A1(n4744), .B0(n4743), .B1(n4414), .C0(n4742), 
        .Y(n4745) );
  OAI221X2 U23 ( .A0(n4416), .A1(n4775), .B0(n4774), .B1(n4414), .C0(n4773), 
        .Y(n4776) );
  OAI221X2 U24 ( .A0(n4416), .A1(n4907), .B0(n4906), .B1(n4413), .C0(n4905), 
        .Y(n4908) );
  OAI221X4 U25 ( .A0(n4416), .A1(n4784), .B0(n4783), .B1(n4413), .C0(n4782), 
        .Y(n4785) );
  OAI221X4 U26 ( .A0(n4415), .A1(n4916), .B0(n4915), .B1(n4413), .C0(n4914), 
        .Y(n4917) );
  OAI221X1 U27 ( .A0(n4407), .A1(n4722), .B0(n4717), .B1(n4404), .C0(n4716), 
        .Y(n4724) );
  INVX3 U28 ( .A(next_RData2[2]), .Y(n4936) );
  INVX3 U29 ( .A(next_RData1[2]), .Y(n4932) );
  INVX3 U30 ( .A(next_RData2[20]), .Y(n4752) );
  OAI221X1 U33 ( .A0(n4416), .A1(n4955), .B0(n4954), .B1(n4413), .C0(n4953), 
        .Y(n4956) );
  INVX3 U35 ( .A(next_RData2[1]), .Y(n4970) );
  XNOR2X2 U38 ( .A(n4839), .B(n4838), .Y(n4850) );
  OAI221X1 U43 ( .A0(n4406), .A1(n4695), .B0(n4690), .B1(n4404), .C0(n4689), 
        .Y(n4697) );
  OAI221X1 U44 ( .A0(n4407), .A1(n4713), .B0(n4708), .B1(n4404), .C0(n4707), 
        .Y(n4715) );
  OAI221X1 U45 ( .A0(n4407), .A1(n4704), .B0(n4699), .B1(n4404), .C0(n4698), 
        .Y(n4706) );
  XNOR2X1 U46 ( .A(n4675), .B(n4674), .Y(n4686) );
  XNOR2X1 U48 ( .A(n4684), .B(n4683), .Y(n4685) );
  OAI221X1 U49 ( .A0(n4407), .A1(n4682), .B0(n4677), .B1(n4404), .C0(n4676), 
        .Y(n4684) );
  NOR2X1 U50 ( .A(n4269), .B(\regfile[1][10] ), .Y(n4204) );
  NAND2X1 U51 ( .A(n4251), .B(n4250), .Y(n3856) );
  MXI2X2 U52 ( .A(n193), .B(n194), .S0(N21), .Y(N138) );
  MXI2X2 U53 ( .A(n226), .B(n227), .S0(n3732), .Y(N122) );
  CLKMX2X2 U54 ( .A(N160), .B(RData2[19]), .S0(n4438), .Y(next_RData2[19]) );
  CLKMX2X2 U55 ( .A(N149), .B(RData2[30]), .S0(n4440), .Y(next_RData2[30]) );
  CLKMX2X2 U56 ( .A(N117), .B(RData1[30]), .S0(n4440), .Y(next_RData1[30]) );
  CLKMX2X2 U57 ( .A(N169), .B(RData2[10]), .S0(n4438), .Y(next_RData2[10]) );
  CLKMX2X2 U58 ( .A(N176), .B(RData2[3]), .S0(n4439), .Y(next_RData2[3]) );
  CLKMX2X2 U59 ( .A(N173), .B(RData2[6]), .S0(n4439), .Y(next_RData2[6]) );
  CLKMX2X2 U60 ( .A(N172), .B(RData2[7]), .S0(n4439), .Y(next_RData2[7]) );
  CLKMX2X2 U61 ( .A(N174), .B(RData2[5]), .S0(n4439), .Y(next_RData2[5]) );
  CLKMX2X2 U62 ( .A(N165), .B(RData2[14]), .S0(n4438), .Y(next_RData2[14]) );
  CLKMX2X2 U63 ( .A(N175), .B(RData2[4]), .S0(n4439), .Y(next_RData2[4]) );
  MX4XL U64 ( .A(n331), .B(n329), .C(n330), .D(n328), .S0(N20), .S1(n3739), 
        .Y(n198) );
  NAND2X2 U65 ( .A(n4246), .B(n4245), .Y(n3864) );
  INVXL U66 ( .A(N18), .Y(n4431) );
  NOR4XL U67 ( .A(N18), .B(n4429), .C(Instruction[9]), .D(Instruction[8]), .Y(
        n185) );
  MXI4XL U68 ( .A(\regfile[8][8] ), .B(\regfile[9][8] ), .C(\regfile[10][8] ), 
        .D(\regfile[11][8] ), .S0(n3769), .S1(N18), .Y(n309) );
  MXI4XL U69 ( .A(\regfile[8][7] ), .B(\regfile[9][7] ), .C(\regfile[10][7] ), 
        .D(\regfile[11][7] ), .S0(n3769), .S1(N18), .Y(n301) );
  MXI4XL U70 ( .A(\regfile[4][7] ), .B(\regfile[5][7] ), .C(\regfile[6][7] ), 
        .D(\regfile[7][7] ), .S0(n3769), .S1(N18), .Y(n302) );
  MXI4XL U71 ( .A(\regfile[12][7] ), .B(\regfile[13][7] ), .C(\regfile[14][7] ), .D(\regfile[15][7] ), .S0(n3768), .S1(N18), .Y(n300) );
  MXI4XL U72 ( .A(\regfile[16][7] ), .B(\regfile[17][7] ), .C(\regfile[18][7] ), .D(\regfile[19][7] ), .S0(n3768), .S1(N18), .Y(n299) );
  MXI4XL U73 ( .A(\regfile[8][6] ), .B(\regfile[9][6] ), .C(\regfile[10][6] ), 
        .D(\regfile[11][6] ), .S0(n3768), .S1(N18), .Y(n293) );
  MXI4XL U74 ( .A(\regfile[24][6] ), .B(\regfile[25][6] ), .C(\regfile[26][6] ), .D(\regfile[27][6] ), .S0(n3768), .S1(N18), .Y(n289) );
  MXI4XL U75 ( .A(\regfile[12][6] ), .B(\regfile[13][6] ), .C(\regfile[14][6] ), .D(\regfile[15][6] ), .S0(n3768), .S1(N18), .Y(n292) );
  MXI4XL U76 ( .A(\regfile[16][6] ), .B(\regfile[17][6] ), .C(\regfile[18][6] ), .D(\regfile[19][6] ), .S0(n3768), .S1(N18), .Y(n291) );
  MXI4XL U77 ( .A(\regfile[4][6] ), .B(\regfile[5][6] ), .C(\regfile[6][6] ), 
        .D(\regfile[7][6] ), .S0(n3768), .S1(N18), .Y(n294) );
  CLKBUFX2 U78 ( .A(N18), .Y(n3741) );
  NAND2X1 U79 ( .A(n4417), .B(MEM_RegWrite), .Y(n4643) );
  MX4X2 U80 ( .A(n327), .B(n325), .C(n326), .D(n324), .S0(N20), .S1(n3739), 
        .Y(n195) );
  MX4X1 U81 ( .A(n319), .B(n317), .C(n318), .D(n316), .S0(N20), .S1(n3739), 
        .Y(n193) );
  MX4X1 U82 ( .A(n351), .B(n349), .C(n350), .D(n348), .S0(N20), .S1(n3739), 
        .Y(n201) );
  MX4X1 U83 ( .A(n311), .B(n309), .C(n310), .D(n308), .S0(N20), .S1(n3739), 
        .Y(n189) );
  MX4X1 U84 ( .A(n447), .B(n445), .C(n446), .D(n444), .S0(n3736), .S1(N19), 
        .Y(n226) );
  MX4X1 U85 ( .A(n439), .B(n437), .C(n438), .D(n436), .S0(n3736), .S1(N19), 
        .Y(n223) );
  MX4X1 U86 ( .A(n431), .B(n429), .C(n430), .D(n428), .S0(n3736), .S1(n3738), 
        .Y(n221) );
  MX4X2 U87 ( .A(n415), .B(n413), .C(n414), .D(n412), .S0(n3736), .S1(N19), 
        .Y(n217) );
  CLKMX2X2 U129 ( .A(N150), .B(RData2[29]), .S0(n4440), .Y(next_RData2[29]) );
  MXI2X2 U130 ( .A(n3835), .B(n3836), .S0(n4257), .Y(N150) );
  CLKMX2X2 U131 ( .A(N155), .B(RData2[24]), .S0(n4440), .Y(next_RData2[24]) );
  MXI2X2 U132 ( .A(n3825), .B(n3826), .S0(n4257), .Y(N155) );
  CLKMX2X2 U133 ( .A(N166), .B(RData2[13]), .S0(n4438), .Y(next_RData2[13]) );
  MXI2X2 U134 ( .A(n3803), .B(n3804), .S0(N26), .Y(N166) );
  CLKMX2X2 U135 ( .A(N154), .B(RData2[25]), .S0(n4440), .Y(next_RData2[25]) );
  MXI2X2 U136 ( .A(n3827), .B(n3828), .S0(n4257), .Y(N154) );
  MXI2X2 U137 ( .A(n1575), .B(n3702), .S0(n3773), .Y(n3705) );
  MXI2X2 U138 ( .A(n236), .B(n237), .S0(n3732), .Y(N117) );
  MXI2X2 U139 ( .A(n203), .B(n204), .S0(N21), .Y(N133) );
  CLKMX2X2 U140 ( .A(N168), .B(RData2[11]), .S0(n4438), .Y(next_RData2[11]) );
  MXI2X2 U141 ( .A(n3799), .B(n3800), .S0(N26), .Y(N168) );
  CLKMX2X2 U142 ( .A(N177), .B(RData2[2]), .S0(n4439), .Y(next_RData2[2]) );
  MXI2X2 U143 ( .A(n3781), .B(n3782), .S0(N26), .Y(N177) );
  CLKMX2X2 U144 ( .A(N171), .B(RData2[8]), .S0(n4438), .Y(next_RData2[8]) );
  MXI2X2 U145 ( .A(n3793), .B(n3794), .S0(N26), .Y(N171) );
  XOR2X2 U146 ( .A(n4861), .B(n4860), .Y(n100) );
  OAI221X2 U147 ( .A0(n4416), .A1(n4859), .B0(n4858), .B1(n4413), .C0(n4857), 
        .Y(n4860) );
  XNOR2X2 U148 ( .A(n4764), .B(n4763), .Y(n4765) );
  CLKMX2X2 U149 ( .A(N170), .B(RData2[9]), .S0(n4438), .Y(next_RData2[9]) );
  MXI2X2 U150 ( .A(n3795), .B(n3796), .S0(N26), .Y(N170) );
  MXI2X2 U151 ( .A(n238), .B(n239), .S0(n3732), .Y(N116) );
  MX4X2 U152 ( .A(n367), .B(n365), .C(n366), .D(n364), .S0(n3735), .S1(N19), 
        .Y(n205) );
  MX4X2 U153 ( .A(n4024), .B(n4022), .C(n4023), .D(n4021), .S0(n4261), .S1(
        n4264), .Y(n3821) );
  MX4X2 U154 ( .A(n3984), .B(n3982), .C(n3983), .D(n3981), .S0(N25), .S1(n4263), .Y(n3811) );
  MXI2X2 U155 ( .A(n3783), .B(n3784), .S0(N26), .Y(N176) );
  MXI2X2 U156 ( .A(n173), .B(n174), .S0(N21), .Y(N141) );
  MXI2X2 U157 ( .A(n160), .B(n161), .S0(N21), .Y(N145) );
  MXI2X2 U158 ( .A(n228), .B(n229), .S0(n3732), .Y(N121) );
  MXI2X2 U159 ( .A(n3787), .B(n3788), .S0(N26), .Y(N174) );
  MXI2X2 U160 ( .A(n175), .B(n188), .S0(N21), .Y(N140) );
  MXI2X2 U161 ( .A(n213), .B(n214), .S0(N21), .Y(N128) );
  MXI2X2 U162 ( .A(n207), .B(n208), .S0(N21), .Y(N131) );
  MXI2X2 U163 ( .A(n164), .B(n165), .S0(N21), .Y(N143) );
  MXI2X2 U164 ( .A(n3823), .B(n3824), .S0(n4257), .Y(N156) );
  MXI2X2 U165 ( .A(n219), .B(n220), .S0(n3732), .Y(N125) );
  MXI2X2 U166 ( .A(n156), .B(n157), .S0(N21), .Y(N147) );
  MXI2X2 U167 ( .A(n3813), .B(n3814), .S0(N26), .Y(N161) );
  MXI2X2 U168 ( .A(n162), .B(n163), .S0(N21), .Y(N144) );
  MXI2X2 U169 ( .A(n3791), .B(n3792), .S0(N26), .Y(N172) );
  MX4X2 U170 ( .A(n3904), .B(n3902), .C(n3903), .D(n3901), .S0(n4259), .S1(
        n4262), .Y(n3791) );
  MXI2X2 U171 ( .A(n3815), .B(n3816), .S0(N26), .Y(N160) );
  MX4X2 U172 ( .A(n4000), .B(n3998), .C(n3999), .D(n3997), .S0(N25), .S1(n4263), .Y(n3815) );
  OAI221X2 U173 ( .A0(n4407), .A1(n4859), .B0(n4854), .B1(n4405), .C0(n4853), 
        .Y(n4861) );
  MX4X2 U175 ( .A(n3896), .B(n3894), .C(n3895), .D(n3893), .S0(n4259), .S1(
        n4262), .Y(n3789) );
  MXI2X2 U176 ( .A(n232), .B(n233), .S0(n3732), .Y(N119) );
  MX4X2 U177 ( .A(n471), .B(n469), .C(n470), .D(n468), .S0(n3737), .S1(n3740), 
        .Y(n232) );
  MXI2X2 U178 ( .A(n230), .B(n231), .S0(n3732), .Y(N120) );
  MX4X2 U179 ( .A(n463), .B(n461), .C(n462), .D(n460), .S0(n3737), .S1(n3740), 
        .Y(n230) );
  MXI2X2 U180 ( .A(n3809), .B(n3810), .S0(N26), .Y(N163) );
  MX4X2 U181 ( .A(n3976), .B(n3974), .C(n3975), .D(n3973), .S0(N25), .S1(n4263), .Y(n3809) );
  MXI2X4 U182 ( .A(n197), .B(n198), .S0(N21), .Y(N136) );
  MXI2X4 U183 ( .A(n199), .B(n200), .S0(N21), .Y(N135) );
  XNOR2X4 U184 ( .A(n4657), .B(n4656), .Y(n4688) );
  OAI221X2 U185 ( .A0(n4415), .A1(n4655), .B0(n4654), .B1(n4414), .C0(n4653), 
        .Y(n4656) );
  MXI2X2 U186 ( .A(n3785), .B(n3786), .S0(N26), .Y(N175) );
  MX4X2 U187 ( .A(n3880), .B(n3878), .C(n3879), .D(n3877), .S0(n4259), .S1(
        n4262), .Y(n3785) );
  MXI2X2 U188 ( .A(n223), .B(n225), .S0(n3732), .Y(N123) );
  MXI2X2 U189 ( .A(n3777), .B(n3778), .S0(n4257), .Y(N179) );
  MX4X2 U190 ( .A(n3848), .B(n3846), .C(n3847), .D(n3845), .S0(N25), .S1(n4264), .Y(n3777) );
  MXI2X2 U191 ( .A(n234), .B(n235), .S0(n3732), .Y(N118) );
  MX4X2 U192 ( .A(n479), .B(n477), .C(n478), .D(n476), .S0(n3737), .S1(n3740), 
        .Y(n234) );
  MXI2X2 U193 ( .A(n201), .B(n202), .S0(N21), .Y(N134) );
  MXI2X2 U194 ( .A(n189), .B(n190), .S0(N21), .Y(N139) );
  XNOR2X4 U195 ( .A(n4821), .B(n4820), .Y(n4852) );
  OAI221X2 U196 ( .A0(n4416), .A1(n4819), .B0(n4818), .B1(n4413), .C0(n4817), 
        .Y(n4820) );
  MXI2X2 U197 ( .A(n209), .B(n210), .S0(N21), .Y(N130) );
  MX4X4 U198 ( .A(n383), .B(n381), .C(n382), .D(n380), .S0(n3735), .S1(N19), 
        .Y(n209) );
  XNOR2X4 U199 ( .A(n4666), .B(n4665), .Y(n4687) );
  OAI221X2 U200 ( .A0(n4415), .A1(n4664), .B0(n4663), .B1(n4414), .C0(n4662), 
        .Y(n4665) );
  NOR2BX2 U201 ( .AN(n4277), .B(\regfile[3][6] ), .Y(n4222) );
  OAI221X4 U202 ( .A0(n4406), .A1(n4655), .B0(n4648), .B1(n4404), .C0(n4647), 
        .Y(n4657) );
  OAI221X2 U203 ( .A0(n4415), .A1(n4673), .B0(n4672), .B1(n4414), .C0(n4671), 
        .Y(n4674) );
  OAI221X2 U204 ( .A0(n4416), .A1(n4837), .B0(n4836), .B1(n4969), .C0(n4835), 
        .Y(n4838) );
  XNOR2X4 U205 ( .A(n4909), .B(n4908), .Y(n4930) );
  OAI221X2 U206 ( .A0(n4415), .A1(n4682), .B0(n4681), .B1(n4414), .C0(n4680), 
        .Y(n4683) );
  OAI221X4 U207 ( .A0(n4963), .A1(n4664), .B0(n4659), .B1(n4961), .C0(n4658), 
        .Y(n4666) );
  XNOR2X4 U208 ( .A(n4715), .B(n4714), .Y(n4726) );
  OAI221X2 U209 ( .A0(n4415), .A1(n4713), .B0(n4712), .B1(n4414), .C0(n4711), 
        .Y(n4714) );
  OAI221X2 U210 ( .A0(n4416), .A1(n4846), .B0(n4845), .B1(n4969), .C0(n4844), 
        .Y(n4847) );
  XNOR2X4 U211 ( .A(n4870), .B(n4869), .Y(n4891) );
  OAI221X2 U212 ( .A0(n4416), .A1(n4868), .B0(n4867), .B1(n4969), .C0(n4866), 
        .Y(n4869) );
  OAI221X2 U213 ( .A0(n4416), .A1(n4877), .B0(n4876), .B1(n4414), .C0(n4875), 
        .Y(n4878) );
  XNOR2X4 U214 ( .A(n4724), .B(n4723), .Y(n4725) );
  OAI221X2 U215 ( .A0(n4415), .A1(n4722), .B0(n4721), .B1(n4414), .C0(n4720), 
        .Y(n4723) );
  XNOR2X4 U216 ( .A(n4888), .B(n4887), .Y(n4889) );
  OAI221X2 U217 ( .A0(n4416), .A1(n4886), .B0(n4885), .B1(n4413), .C0(n4884), 
        .Y(n4887) );
  XNOR2X4 U218 ( .A(n4786), .B(n4785), .Y(n4807) );
  XNOR2X4 U219 ( .A(n4918), .B(n4917), .Y(n4929) );
  XNOR2X4 U220 ( .A(n4804), .B(n4803), .Y(n4805) );
  OAI221X2 U221 ( .A0(n4416), .A1(n4802), .B0(n4801), .B1(n4414), .C0(n4800), 
        .Y(n4803) );
  OAI221X2 U222 ( .A0(n4416), .A1(n4971), .B0(n4970), .B1(n4413), .C0(n4968), 
        .Y(n4973) );
  MXI2X4 U223 ( .A(n158), .B(n159), .S0(N21), .Y(N146) );
  MX4X4 U224 ( .A(n255), .B(n253), .C(n254), .D(n252), .S0(n3733), .S1(n3740), 
        .Y(n158) );
  OAI221X2 U225 ( .A0(n4415), .A1(n4753), .B0(n4752), .B1(n4414), .C0(n4751), 
        .Y(n4754) );
  XNOR2X4 U226 ( .A(n4927), .B(n4926), .Y(n4928) );
  OAI221X2 U227 ( .A0(n4416), .A1(n4925), .B0(n4924), .B1(n4413), .C0(n4923), 
        .Y(n4926) );
  OAI221X2 U228 ( .A0(n4415), .A1(n4762), .B0(n4761), .B1(n4414), .C0(n4760), 
        .Y(n4763) );
  INVX4 U229 ( .A(next_RData2[21]), .Y(n4761) );
  MXI2X2 U230 ( .A(n1579), .B(n4247), .S0(n4297), .Y(n4250) );
  OAI221X4 U231 ( .A0(n4406), .A1(n4886), .B0(n4881), .B1(n4405), .C0(n4880), 
        .Y(n4888) );
  XNOR2X4 U232 ( .A(n4777), .B(n4776), .Y(n4808) );
  OAI221X1 U233 ( .A0(n4407), .A1(n4775), .B0(n4770), .B1(n4405), .C0(n4769), 
        .Y(n4777) );
  NOR2X6 U234 ( .A(n4204), .B(n4203), .Y(n4206) );
  XNOR2X4 U235 ( .A(n4746), .B(n4745), .Y(n4767) );
  OAI221X2 U237 ( .A0(n4406), .A1(n4925), .B0(n4920), .B1(n4961), .C0(n4919), 
        .Y(n4927) );
  NAND2X2 U238 ( .A(n3726), .B(n3725), .Y(n255) );
  MXI2X2 U239 ( .A(n1579), .B(n3722), .S0(n3772), .Y(n3725) );
  XNOR2X1 U240 ( .A(n4755), .B(n4754), .Y(n4766) );
  XNOR2X4 U243 ( .A(n4697), .B(n4696), .Y(n4728) );
  OAI221X2 U244 ( .A0(n4415), .A1(n4695), .B0(n4694), .B1(n4414), .C0(n4693), 
        .Y(n4696) );
  XNOR2X4 U245 ( .A(n4830), .B(n4829), .Y(n4851) );
  OAI221X2 U246 ( .A0(n4416), .A1(n4828), .B0(n4827), .B1(n4413), .C0(n4826), 
        .Y(n4829) );
  XNOR2X4 U247 ( .A(n4706), .B(n4705), .Y(n4727) );
  OAI221X2 U248 ( .A0(n4415), .A1(n4704), .B0(n4703), .B1(n4414), .C0(n4702), 
        .Y(n4705) );
  OAI221X2 U250 ( .A0(n4415), .A1(n4898), .B0(n4897), .B1(n4413), .C0(n4896), 
        .Y(n4899) );
  XNOR2X4 U251 ( .A(n4737), .B(n4736), .Y(n4768) );
  OAI221X2 U252 ( .A0(n4415), .A1(n4735), .B0(n4734), .B1(n4414), .C0(n4733), 
        .Y(n4736) );
  OAI221X2 U253 ( .A0(n4415), .A1(n4937), .B0(n4936), .B1(n4413), .C0(n4935), 
        .Y(n4938) );
  MXI2X4 U254 ( .A(n217), .B(n218), .S0(n3732), .Y(N126) );
  MXI2X4 U255 ( .A(n215), .B(n216), .S0(n3732), .Y(N127) );
  MX4X4 U256 ( .A(n407), .B(n405), .C(n406), .D(n404), .S0(n3736), .S1(n3739), 
        .Y(n215) );
  MXI2X4 U257 ( .A(n221), .B(n222), .S0(n3732), .Y(N124) );
  MXI2X4 U258 ( .A(n195), .B(n196), .S0(N21), .Y(N137) );
  MXI2X4 U259 ( .A(n211), .B(n212), .S0(N21), .Y(N129) );
  MX4X4 U260 ( .A(n391), .B(n389), .C(n390), .D(n388), .S0(n3735), .S1(N19), 
        .Y(n211) );
  CLKAND2X6 U261 ( .A(n4269), .B(n1545), .Y(n4237) );
  XNOR2X4 U262 ( .A(n4948), .B(n4947), .Y(n4977) );
  OAI221X2 U263 ( .A0(n4972), .A1(n4946), .B0(n4945), .B1(n4413), .C0(n4944), 
        .Y(n4947) );
  NOR2X6 U264 ( .A(n102), .B(n103), .Y(equal) );
  OR4X6 U265 ( .A(n4981), .B(n4980), .C(n4979), .D(n4978), .Y(n103) );
  OR4X6 U266 ( .A(n4812), .B(n4811), .C(n4810), .D(n4809), .Y(n102) );
  OAI221X2 U267 ( .A0(n4406), .A1(n4937), .B0(n4932), .B1(n4405), .C0(n4931), 
        .Y(n4939) );
  OR2X4 U269 ( .A(n4893), .B(n4961), .Y(n96) );
  OR2XL U270 ( .A(n4406), .B(n4898), .Y(n95) );
  NOR2X1 U272 ( .A(\regfile[1][6] ), .B(n4275), .Y(n4224) );
  NOR2X1 U273 ( .A(\regfile[1][2] ), .B(n4275), .Y(n4244) );
  XOR2X1 U274 ( .A(n4938), .B(n4939), .Y(n99) );
  INVX3 U275 ( .A(EX_RegWriteData[30]), .Y(n4655) );
  INVXL U276 ( .A(N24), .Y(n4425) );
  INVXL U277 ( .A(N20), .Y(n4434) );
  INVXL U278 ( .A(N19), .Y(n4432) );
  NOR2X1 U281 ( .A(n4275), .B(\regfile[1][7] ), .Y(n4219) );
  NOR2X1 U285 ( .A(n4278), .B(\regfile[1][16] ), .Y(n4174) );
  NOR2X1 U286 ( .A(n4276), .B(\regfile[1][17] ), .Y(n4169) );
  NOR2X1 U287 ( .A(n4280), .B(\regfile[1][18] ), .Y(n4164) );
  NOR2X1 U289 ( .A(n4277), .B(\regfile[1][20] ), .Y(n4154) );
  NOR2X1 U290 ( .A(n4269), .B(\regfile[1][23] ), .Y(n4139) );
  NOR2X1 U291 ( .A(n4268), .B(\regfile[1][21] ), .Y(n4149) );
  NOR2X1 U292 ( .A(n4270), .B(\regfile[1][22] ), .Y(n4144) );
  NOR2X1 U294 ( .A(n4277), .B(\regfile[1][27] ), .Y(n4119) );
  NOR2X1 U295 ( .A(\regfile[1][25] ), .B(n4274), .Y(n4129) );
  NOR2X1 U296 ( .A(n4270), .B(\regfile[1][26] ), .Y(n4124) );
  NOR2X1 U297 ( .A(n4268), .B(\regfile[1][15] ), .Y(n4179) );
  NOR2X1 U298 ( .A(n4277), .B(\regfile[1][31] ), .Y(n4099) );
  NOR2X1 U299 ( .A(n4275), .B(\regfile[1][28] ), .Y(n4114) );
  NOR2X1 U300 ( .A(\regfile[1][29] ), .B(n4279), .Y(n4109) );
  NOR2X1 U301 ( .A(n4270), .B(\regfile[1][30] ), .Y(n4104) );
  NOR2X1 U302 ( .A(\regfile[1][8] ), .B(n4270), .Y(n4214) );
  NOR2X1 U304 ( .A(n4280), .B(\regfile[1][12] ), .Y(n4194) );
  NOR2X1 U305 ( .A(n4274), .B(\regfile[1][13] ), .Y(n4189) );
  NOR2X1 U306 ( .A(n4276), .B(\regfile[1][14] ), .Y(n4184) );
  NOR2X1 U307 ( .A(\regfile[1][1] ), .B(n4274), .Y(n4249) );
  NOR2BX1 U308 ( .AN(n4276), .B(n94), .Y(n4157) );
  NOR2BX1 U309 ( .AN(n4279), .B(\regfile[3][16] ), .Y(n4172) );
  NOR2BX1 U310 ( .AN(n4269), .B(\regfile[3][17] ), .Y(n4167) );
  NOR2BX1 U311 ( .AN(n4274), .B(n91), .Y(n4162) );
  NOR2BX1 U312 ( .AN(n4268), .B(n85), .Y(n4152) );
  NOR2BX1 U313 ( .AN(n4268), .B(n87), .Y(n4137) );
  NOR2BX1 U314 ( .AN(n4268), .B(\regfile[3][21] ), .Y(n4147) );
  NOR2BX1 U315 ( .AN(n4278), .B(n89), .Y(n4217) );
  NOR2BX1 U316 ( .AN(n4268), .B(\regfile[3][22] ), .Y(n4142) );
  NOR2BX1 U317 ( .AN(n4268), .B(\regfile[3][9] ), .Y(n4207) );
  NOR2BX1 U318 ( .AN(n4274), .B(\regfile[3][8] ), .Y(n4212) );
  NOR2BX1 U319 ( .AN(n4277), .B(\regfile[3][11] ), .Y(n4197) );
  NOR2BX1 U320 ( .AN(n4276), .B(\regfile[3][24] ), .Y(n4132) );
  NOR2BX1 U321 ( .AN(n4270), .B(\regfile[3][15] ), .Y(n4177) );
  NOR2BX1 U322 ( .AN(n4275), .B(\regfile[3][13] ), .Y(n4187) );
  NOR2BX1 U323 ( .AN(n4277), .B(\regfile[3][14] ), .Y(n4182) );
  NOR2BX1 U324 ( .AN(n4269), .B(\regfile[3][5] ), .Y(n4227) );
  NOR2BX1 U325 ( .AN(n4280), .B(n92), .Y(n4252) );
  NOR2BX1 U326 ( .AN(n4278), .B(\regfile[3][2] ), .Y(n4242) );
  NOR2BX1 U327 ( .AN(n4269), .B(n90), .Y(n4232) );
  NOR2BX1 U328 ( .AN(n4269), .B(\regfile[3][27] ), .Y(n4117) );
  NOR2BX1 U329 ( .AN(n4275), .B(\regfile[3][25] ), .Y(n4127) );
  NOR2BX1 U330 ( .AN(n4279), .B(\regfile[3][26] ), .Y(n4122) );
  NOR2BX1 U331 ( .AN(n4274), .B(\regfile[3][12] ), .Y(n4192) );
  NOR2BX1 U332 ( .AN(n4280), .B(\regfile[3][31] ), .Y(n4097) );
  NOR2BX1 U333 ( .AN(n4268), .B(\regfile[3][28] ), .Y(n4112) );
  NOR2BX1 U334 ( .AN(n4269), .B(\regfile[3][29] ), .Y(n4107) );
  NOR2BX1 U335 ( .AN(n4270), .B(\regfile[3][30] ), .Y(n4102) );
  NOR2BX1 U336 ( .AN(n4270), .B(\regfile[3][1] ), .Y(n4247) );
  NAND4X2 U337 ( .A(n4728), .B(n4727), .C(n4726), .D(n4725), .Y(n4811) );
  NAND2X2 U338 ( .A(Branch), .B(equal), .Y(n4982) );
  NAND4X2 U339 ( .A(n4768), .B(n4767), .C(n4766), .D(n4765), .Y(n4810) );
  NAND4X2 U340 ( .A(n4808), .B(n4807), .C(n4806), .D(n4805), .Y(n4809) );
  NAND4X2 U341 ( .A(n4685), .B(n4687), .C(n4686), .D(n4688), .Y(n4812) );
  NAND4X2 U342 ( .A(n4852), .B(n4851), .C(n4850), .D(n4849), .Y(n4981) );
  NAND4BX2 U344 ( .AN(n99), .B(n4977), .C(n4976), .D(n4975), .Y(n4978) );
  NAND4BX2 U345 ( .AN(n100), .B(n4891), .C(n4890), .D(n4889), .Y(n4980) );
  CLKINVX1 U346 ( .A(n4423), .Y(n4422) );
  CLKINVX1 U347 ( .A(stall), .Y(n4448) );
  CLKINVX1 U348 ( .A(N22), .Y(n4423) );
  CLKINVX1 U349 ( .A(N25), .Y(n4427) );
  CLKINVX1 U350 ( .A(N17), .Y(n4430) );
  CLKINVX1 U351 ( .A(N23), .Y(n4424) );
  CLKINVX1 U352 ( .A(N26), .Y(n4428) );
  CLKINVX1 U353 ( .A(N21), .Y(n4435) );
  CLKMX2X4 U354 ( .A(N151), .B(RData2[28]), .S0(n4439), .Y(next_RData2[28]) );
  CLKMX2X4 U355 ( .A(N116), .B(RData1[31]), .S0(n4440), .Y(next_RData1[31]) );
  CLKMX2X4 U356 ( .A(N121), .B(RData1[26]), .S0(n4440), .Y(next_RData1[26]) );
  CLKMX2X4 U357 ( .A(N120), .B(RData1[27]), .S0(n4440), .Y(next_RData1[27]) );
  CLKMX2X4 U358 ( .A(N119), .B(RData1[28]), .S0(n4439), .Y(next_RData1[28]) );
  CLKMX2X4 U359 ( .A(N122), .B(RData1[25]), .S0(n4440), .Y(next_RData1[25]) );
  CLKMX2X4 U360 ( .A(N118), .B(RData1[29]), .S0(n4439), .Y(next_RData1[29]) );
  CLKMX2X4 U361 ( .A(N128), .B(RData1[19]), .S0(n4437), .Y(next_RData1[19]) );
  CLKMX2X4 U362 ( .A(N125), .B(RData1[22]), .S0(n4440), .Y(next_RData1[22]) );
  CLKMX2X4 U363 ( .A(N145), .B(RData1[2]), .S0(n4439), .Y(next_RData1[2]) );
  CLKMX2X4 U364 ( .A(N147), .B(RData1[0]), .S0(n4439), .Y(next_RData1[0]) );
  CLKMX2X4 U365 ( .A(N127), .B(RData1[20]), .S0(n4440), .Y(next_RData1[20]) );
  CLKMX2X4 U366 ( .A(N144), .B(RData1[3]), .S0(n4439), .Y(next_RData1[3]) );
  CLKMX2X4 U367 ( .A(N123), .B(RData1[24]), .S0(n4440), .Y(next_RData1[24]) );
  CLKMX2X4 U368 ( .A(N143), .B(RData1[4]), .S0(n4439), .Y(next_RData1[4]) );
  CLKMX2X4 U369 ( .A(N141), .B(RData1[6]), .S0(n4439), .Y(next_RData1[6]) );
  CLKMX2X4 U370 ( .A(N140), .B(RData1[7]), .S0(n4439), .Y(next_RData1[7]) );
  CLKMX2X4 U371 ( .A(N126), .B(RData1[21]), .S0(n4440), .Y(next_RData1[21]) );
  CLKMX2X4 U372 ( .A(N146), .B(RData1[1]), .S0(n4439), .Y(next_RData1[1]) );
  CLKMX2X4 U373 ( .A(N142), .B(RData1[5]), .S0(n4439), .Y(next_RData1[5]) );
  CLKMX2X4 U374 ( .A(N132), .B(RData1[15]), .S0(n4438), .Y(next_RData1[15]) );
  CLKMX2X4 U375 ( .A(N133), .B(RData1[14]), .S0(n4438), .Y(next_RData1[14]) );
  CLKMX2X4 U376 ( .A(N136), .B(RData1[11]), .S0(n4438), .Y(next_RData1[11]) );
  CLKMX2X4 U377 ( .A(N137), .B(RData1[10]), .S0(n4438), .Y(next_RData1[10]) );
  CLKMX2X4 U378 ( .A(N135), .B(RData1[12]), .S0(n4438), .Y(next_RData1[12]) );
  CLKMX2X4 U379 ( .A(N139), .B(RData1[8]), .S0(n4438), .Y(next_RData1[8]) );
  CLKMX2X4 U380 ( .A(N138), .B(RData1[9]), .S0(n4438), .Y(next_RData1[9]) );
  CLKMX2X4 U381 ( .A(N134), .B(RData1[13]), .S0(n4438), .Y(next_RData1[13]) );
  CLKMX2X4 U382 ( .A(N124), .B(RData1[23]), .S0(n4441), .Y(next_RData1[23]) );
  CLKMX2X4 U383 ( .A(N129), .B(RData1[18]), .S0(n4441), .Y(next_RData1[18]) );
  CLKMX2X4 U384 ( .A(N131), .B(RData1[16]), .S0(n4441), .Y(next_RData1[16]) );
  CLKMX2X4 U385 ( .A(N130), .B(RData1[17]), .S0(n4441), .Y(next_RData1[17]) );
  INVXL U386 ( .A(BranchTaken), .Y(n4989) );
  CLKMX2X4 U387 ( .A(N148), .B(RData2[31]), .S0(n4440), .Y(next_RData2[31]) );
  CLKMX2X4 U388 ( .A(N157), .B(RData2[22]), .S0(n4440), .Y(next_RData2[22]) );
  CLKMX2X4 U389 ( .A(N179), .B(RData2[0]), .S0(n4439), .Y(next_RData2[0]) );
  CLKMX2X4 U390 ( .A(N159), .B(RData2[20]), .S0(n4440), .Y(next_RData2[20]) );
  CLKMX2X4 U391 ( .A(N153), .B(RData2[26]), .S0(n4440), .Y(next_RData2[26]) );
  CLKMX2X4 U392 ( .A(N152), .B(RData2[27]), .S0(n4440), .Y(next_RData2[27]) );
  CLKMX2X4 U393 ( .A(N158), .B(RData2[21]), .S0(n4440), .Y(next_RData2[21]) );
  CLKMX2X4 U394 ( .A(N178), .B(RData2[1]), .S0(n4439), .Y(next_RData2[1]) );
  CLKMX2X4 U395 ( .A(N164), .B(RData2[15]), .S0(n4438), .Y(next_RData2[15]) );
  CLKMX2X4 U396 ( .A(N167), .B(RData2[12]), .S0(n4438), .Y(next_RData2[12]) );
  CLKMX2X4 U397 ( .A(N156), .B(RData2[23]), .S0(n4441), .Y(next_RData2[23]) );
  CLKMX2X4 U398 ( .A(N161), .B(RData2[18]), .S0(n4441), .Y(next_RData2[18]) );
  CLKMX2X4 U399 ( .A(N163), .B(RData2[16]), .S0(n4441), .Y(next_RData2[16]) );
  CLKMX2X4 U400 ( .A(N162), .B(RData2[17]), .S0(n4441), .Y(next_RData2[17]) );
  INVXL U401 ( .A(PCadd4[2]), .Y(n4580) );
  INVXL U402 ( .A(PCadd4[3]), .Y(n4582) );
  INVXL U403 ( .A(PCadd4[4]), .Y(n4584) );
  NAND3XL U404 ( .A(Jump), .B(Instruction[27]), .C(n224), .Y(n191) );
  AND3XL U405 ( .A(Instruction[26]), .B(n4983), .C(n170), .Y(n224) );
  NOR2BXL U406 ( .AN(Reg_W[3]), .B(n4984), .Y(n93) );
  INVX1 U407 ( .A(MEM_RegWrite), .Y(n4983) );
  INVXL U408 ( .A(Reg_W[2]), .Y(n4984) );
  NOR2XL U409 ( .A(Reg_W[2]), .B(Reg_W[3]), .Y(n62) );
  NOR2BXL U410 ( .AN(Reg_W[3]), .B(Reg_W[2]), .Y(n83) );
  NOR2XL U411 ( .A(n4984), .B(Reg_W[3]), .Y(n73) );
  NAND2XL U412 ( .A(Reg_W[1]), .B(Reg_W[0]), .Y(n124) );
  MX2XL U413 ( .A(n4542), .B(WriteData[0]), .S0(n4305), .Y(n1678) );
  MX2XL U414 ( .A(n4543), .B(WriteData[1]), .S0(n4305), .Y(n1680) );
  MX2XL U415 ( .A(n4544), .B(WriteData[2]), .S0(n4305), .Y(n1682) );
  MX2XL U416 ( .A(n4545), .B(WriteData[3]), .S0(n4305), .Y(n1684) );
  MX2XL U417 ( .A(n4546), .B(WriteData[4]), .S0(n4305), .Y(n1686) );
  MX2XL U418 ( .A(n4547), .B(WriteData[5]), .S0(n4305), .Y(n1688) );
  MX2XL U419 ( .A(n4548), .B(WriteData[6]), .S0(n4305), .Y(n1690) );
  MX2XL U420 ( .A(n4549), .B(WriteData[7]), .S0(n4305), .Y(n1692) );
  MX2XL U421 ( .A(n4550), .B(WriteData[8]), .S0(n4305), .Y(n1694) );
  MX2XL U422 ( .A(n4551), .B(WriteData[9]), .S0(n4305), .Y(n1696) );
  MX2XL U423 ( .A(n4552), .B(WriteData[10]), .S0(n4305), .Y(n1698) );
  MX2XL U424 ( .A(n4553), .B(WriteData[11]), .S0(n4305), .Y(n1700) );
  MX2XL U425 ( .A(n4554), .B(WriteData[12]), .S0(n4305), .Y(n1702) );
  MX2XL U426 ( .A(n4555), .B(WriteData[13]), .S0(n4306), .Y(n1704) );
  MX2XL U427 ( .A(n4556), .B(WriteData[14]), .S0(n4306), .Y(n1706) );
  MX2XL U428 ( .A(n4557), .B(WriteData[15]), .S0(n4306), .Y(n1708) );
  MX2XL U429 ( .A(n4558), .B(WriteData[16]), .S0(n4306), .Y(n1710) );
  MX2XL U430 ( .A(n4559), .B(WriteData[17]), .S0(n4306), .Y(n1712) );
  MX2XL U431 ( .A(n4560), .B(WriteData[18]), .S0(n4306), .Y(n1714) );
  MX2XL U432 ( .A(n4561), .B(WriteData[19]), .S0(n4306), .Y(n1716) );
  MX2XL U433 ( .A(n4562), .B(WriteData[20]), .S0(n4306), .Y(n1718) );
  MX2XL U434 ( .A(n4563), .B(WriteData[21]), .S0(n4306), .Y(n1720) );
  MX2XL U435 ( .A(n4564), .B(WriteData[22]), .S0(n4306), .Y(n1722) );
  MX2XL U436 ( .A(n4565), .B(WriteData[23]), .S0(n4306), .Y(n1724) );
  MX2XL U437 ( .A(n4566), .B(WriteData[24]), .S0(n4306), .Y(n1726) );
  MX2XL U438 ( .A(n4567), .B(WriteData[25]), .S0(n4306), .Y(n1728) );
  MX2XL U439 ( .A(n4568), .B(WriteData[26]), .S0(n114), .Y(n1730) );
  MX2XL U440 ( .A(n4569), .B(WriteData[27]), .S0(n4305), .Y(n1732) );
  MX2XL U441 ( .A(n4572), .B(WriteData[30]), .S0(n4306), .Y(n1738) );
  MX2XL U442 ( .A(n4573), .B(WriteData[31]), .S0(n114), .Y(n1740) );
  CLKBUFX3 U443 ( .A(n10), .Y(n4302) );
  AO21XL U444 ( .A0(Instruction[28]), .A1(Instruction[29]), .B0(n12), .Y(n10)
         );
  OAI21XL U445 ( .A0(n613), .A1(n4445), .B0(n4302), .Y(next_Immediate_SE[20])
         );
  OAI21XL U446 ( .A0(n614), .A1(n4445), .B0(n4302), .Y(next_Immediate_SE[21])
         );
  OAI21XL U447 ( .A0(n615), .A1(n4445), .B0(n4302), .Y(next_Immediate_SE[22])
         );
  OAI21XL U448 ( .A0(n616), .A1(n4445), .B0(n4302), .Y(next_Immediate_SE[23])
         );
  OAI21XL U449 ( .A0(n608), .A1(n4445), .B0(n4302), .Y(next_Immediate_SE[16])
         );
  OAI21XL U450 ( .A0(n609), .A1(n4445), .B0(n4302), .Y(next_Immediate_SE[17])
         );
  OAI21XL U451 ( .A0(n610), .A1(n4445), .B0(n4302), .Y(next_Immediate_SE[18])
         );
  OAI21XL U452 ( .A0(n611), .A1(n4445), .B0(n4302), .Y(next_Immediate_SE[19])
         );
  MX2XL U453 ( .A(Instruction[8]), .B(Immediate_SE[8]), .S0(n4437), .Y(n147)
         );
  OAI21XL U454 ( .A0(n617), .A1(n4445), .B0(n4302), .Y(next_Immediate_SE[24])
         );
  OAI21XL U455 ( .A0(n618), .A1(n4445), .B0(n4302), .Y(next_Immediate_SE[25])
         );
  OAI21XL U456 ( .A0(n607), .A1(n4445), .B0(n12), .Y(next_Immediate_SE[15]) );
  MX2XL U457 ( .A(Instruction[6]), .B(Immediate_SE[6]), .S0(n4437), .Y(n149)
         );
  MX2XL U458 ( .A(Instruction[7]), .B(Immediate_SE[7]), .S0(n4437), .Y(n150)
         );
  MX2XL U459 ( .A(Instruction[9]), .B(Immediate_SE[9]), .S0(n4437), .Y(n151)
         );
  MX2XL U460 ( .A(Instruction[2]), .B(n1913), .S0(n4438), .Y(n143) );
  OAI21XL U461 ( .A0(n619), .A1(n4445), .B0(n4302), .Y(next_Immediate_SE[26])
         );
  OAI21XL U462 ( .A0(n620), .A1(n4445), .B0(n4302), .Y(next_Immediate_SE[27])
         );
  OAI21XL U463 ( .A0(n621), .A1(n4445), .B0(n4302), .Y(next_Immediate_SE[28])
         );
  OAI21XL U464 ( .A0(n622), .A1(n4445), .B0(n4302), .Y(next_Immediate_SE[29])
         );
  AND3XL U465 ( .A(Instruction[27]), .B(n170), .C(Instruction[26]), .Y(n169)
         );
  NAND4XL U466 ( .A(Instruction[27]), .B(Instruction[26]), .C(n170), .D(
        MEM_RegWrite), .Y(n167) );
  NOR4XL U467 ( .A(Instruction[4]), .B(Instruction[3]), .C(Instruction[2]), 
        .D(Instruction[27]), .Y(n183) );
  CLKBUFX3 U468 ( .A(n4281), .Y(n4300) );
  CLKBUFX3 U469 ( .A(n4429), .Y(n3775) );
  CLKBUFX3 U470 ( .A(N23), .Y(n4274) );
  CLKBUFX3 U471 ( .A(N18), .Y(n3749) );
  CLKBUFX3 U472 ( .A(n4282), .Y(n4298) );
  CLKBUFX3 U473 ( .A(n4282), .Y(n4299) );
  CLKBUFX3 U474 ( .A(n3757), .Y(n3773) );
  CLKBUFX3 U475 ( .A(n3757), .Y(n3774) );
  CLKBUFX3 U476 ( .A(n4282), .Y(n4297) );
  CLKBUFX3 U477 ( .A(n3756), .Y(n3772) );
  CLKBUFX3 U478 ( .A(n4281), .Y(n4291) );
  CLKBUFX3 U479 ( .A(n4281), .Y(n4292) );
  CLKBUFX3 U480 ( .A(n4282), .Y(n4293) );
  CLKBUFX3 U481 ( .A(n4281), .Y(n4295) );
  CLKBUFX3 U482 ( .A(n4282), .Y(n4296) );
  CLKBUFX3 U483 ( .A(n4281), .Y(n4294) );
  CLKBUFX3 U484 ( .A(n4282), .Y(n4283) );
  CLKBUFX3 U485 ( .A(n4422), .Y(n4284) );
  CLKBUFX3 U486 ( .A(n4281), .Y(n4285) );
  CLKBUFX3 U487 ( .A(n4282), .Y(n4287) );
  CLKBUFX3 U488 ( .A(n4282), .Y(n4288) );
  CLKBUFX3 U489 ( .A(n4281), .Y(n4289) );
  CLKBUFX3 U490 ( .A(n4281), .Y(n4290) );
  CLKBUFX3 U491 ( .A(n4281), .Y(n4286) );
  CLKBUFX3 U492 ( .A(n3756), .Y(n3766) );
  CLKBUFX3 U493 ( .A(n3757), .Y(n3767) );
  CLKBUFX3 U494 ( .A(n3756), .Y(n3768) );
  CLKBUFX3 U495 ( .A(n3756), .Y(n3770) );
  CLKBUFX3 U496 ( .A(n3756), .Y(n3771) );
  CLKBUFX3 U497 ( .A(n3756), .Y(n3769) );
  CLKBUFX3 U498 ( .A(n3757), .Y(n3758) );
  CLKBUFX3 U499 ( .A(n3756), .Y(n3759) );
  CLKBUFX3 U500 ( .A(n3757), .Y(n3760) );
  CLKBUFX3 U501 ( .A(n3757), .Y(n3762) );
  CLKBUFX3 U502 ( .A(n3757), .Y(n3763) );
  CLKBUFX3 U503 ( .A(n3756), .Y(n3764) );
  CLKBUFX3 U504 ( .A(n3756), .Y(n3765) );
  CLKBUFX3 U505 ( .A(n3757), .Y(n3761) );
  BUFX4 U506 ( .A(n4273), .Y(n4271) );
  BUFX4 U507 ( .A(n4266), .Y(n4273) );
  BUFX4 U508 ( .A(n4267), .Y(n4272) );
  BUFX4 U509 ( .A(N23), .Y(n4266) );
  BUFX4 U510 ( .A(N23), .Y(n4267) );
  BUFX4 U511 ( .A(N23), .Y(n4269) );
  BUFX4 U512 ( .A(N23), .Y(n4270) );
  BUFX4 U513 ( .A(N23), .Y(n4268) );
  BUFX4 U514 ( .A(n3741), .Y(n3746) );
  BUFX4 U515 ( .A(n3750), .Y(n3747) );
  BUFX4 U516 ( .A(n3741), .Y(n3748) );
  BUFX4 U517 ( .A(n3741), .Y(n3742) );
  BUFX4 U518 ( .A(n3741), .Y(n3743) );
  BUFX4 U519 ( .A(n3750), .Y(n3744) );
  BUFX4 U520 ( .A(n3750), .Y(n3745) );
  CLKBUFX3 U521 ( .A(N23), .Y(n4275) );
  CLKBUFX3 U522 ( .A(N18), .Y(n3750) );
  CLKBUFX3 U523 ( .A(n4282), .Y(n4301) );
  CLKBUFX3 U524 ( .A(n3757), .Y(n3776) );
  CLKBUFX3 U525 ( .A(N23), .Y(n4276) );
  CLKBUFX3 U526 ( .A(N23), .Y(n4277) );
  CLKBUFX3 U527 ( .A(N23), .Y(n4278) );
  CLKBUFX3 U528 ( .A(N23), .Y(n4279) );
  CLKBUFX3 U529 ( .A(n3741), .Y(n3751) );
  CLKBUFX3 U530 ( .A(n3741), .Y(n3752) );
  CLKBUFX3 U531 ( .A(n3741), .Y(n3753) );
  CLKBUFX3 U532 ( .A(n3741), .Y(n3754) );
  CLKBUFX3 U533 ( .A(n4258), .Y(n4259) );
  CLKBUFX3 U535 ( .A(n4258), .Y(n4261) );
  CLKBUFX3 U536 ( .A(n3733), .Y(n3734) );
  CLKBUFX3 U537 ( .A(n3733), .Y(n3735) );
  CLKBUFX3 U538 ( .A(n3733), .Y(n3736) );
  CLKBUFX3 U539 ( .A(n4433), .Y(n3737) );
  CLKBUFX3 U540 ( .A(N23), .Y(n4280) );
  CLKBUFX3 U541 ( .A(n3741), .Y(n3755) );
  CLKBUFX3 U542 ( .A(N24), .Y(n4262) );
  CLKBUFX3 U543 ( .A(N24), .Y(n4263) );
  CLKBUFX3 U544 ( .A(N24), .Y(n4264) );
  CLKBUFX3 U545 ( .A(N24), .Y(n4265) );
  CLKBUFX3 U546 ( .A(N19), .Y(n3738) );
  CLKBUFX3 U547 ( .A(N19), .Y(n3739) );
  CLKBUFX3 U548 ( .A(N19), .Y(n3740) );
  CLKBUFX3 U549 ( .A(n4969), .Y(n4414) );
  CLKBUFX3 U550 ( .A(n4961), .Y(n4404) );
  CLKBUFX3 U551 ( .A(n4961), .Y(n4405) );
  CLKBUFX3 U552 ( .A(n4422), .Y(n4282) );
  CLKBUFX3 U553 ( .A(n4531), .Y(n4462) );
  CLKBUFX3 U554 ( .A(n4519), .Y(n4513) );
  CLKBUFX3 U555 ( .A(n4519), .Y(n4512) );
  CLKBUFX3 U556 ( .A(n4519), .Y(n4511) );
  CLKBUFX3 U557 ( .A(n4519), .Y(n4510) );
  CLKBUFX3 U558 ( .A(n4520), .Y(n4509) );
  CLKBUFX3 U559 ( .A(n4520), .Y(n4508) );
  CLKBUFX3 U560 ( .A(n4520), .Y(n4507) );
  CLKBUFX3 U561 ( .A(n4520), .Y(n4506) );
  CLKBUFX3 U562 ( .A(n4521), .Y(n4505) );
  CLKBUFX3 U563 ( .A(n4521), .Y(n4504) );
  CLKBUFX3 U564 ( .A(n4521), .Y(n4503) );
  CLKBUFX3 U565 ( .A(n4521), .Y(n4502) );
  CLKBUFX3 U566 ( .A(n4522), .Y(n4501) );
  CLKBUFX3 U567 ( .A(n4522), .Y(n4500) );
  CLKBUFX3 U568 ( .A(n4522), .Y(n4499) );
  CLKBUFX3 U569 ( .A(n4522), .Y(n4498) );
  CLKBUFX3 U570 ( .A(n4523), .Y(n4497) );
  CLKBUFX3 U571 ( .A(n4523), .Y(n4496) );
  CLKBUFX3 U572 ( .A(n4523), .Y(n4495) );
  CLKBUFX3 U573 ( .A(n4523), .Y(n4494) );
  CLKBUFX3 U574 ( .A(n4524), .Y(n4493) );
  CLKBUFX3 U575 ( .A(n4524), .Y(n4492) );
  CLKBUFX3 U576 ( .A(n4524), .Y(n4491) );
  CLKBUFX3 U577 ( .A(n4524), .Y(n4490) );
  CLKBUFX3 U578 ( .A(n4525), .Y(n4489) );
  CLKBUFX3 U579 ( .A(n4525), .Y(n4488) );
  CLKBUFX3 U580 ( .A(n4525), .Y(n4487) );
  CLKBUFX3 U581 ( .A(n4525), .Y(n4486) );
  CLKBUFX3 U582 ( .A(n4526), .Y(n4485) );
  CLKBUFX3 U583 ( .A(n4526), .Y(n4484) );
  CLKBUFX3 U584 ( .A(n4526), .Y(n4483) );
  CLKBUFX3 U585 ( .A(n4526), .Y(n4482) );
  CLKBUFX3 U586 ( .A(n4527), .Y(n4481) );
  CLKBUFX3 U587 ( .A(n4527), .Y(n4480) );
  CLKBUFX3 U588 ( .A(n4527), .Y(n4479) );
  CLKBUFX3 U589 ( .A(n4527), .Y(n4478) );
  CLKBUFX3 U590 ( .A(n4528), .Y(n4477) );
  CLKBUFX3 U591 ( .A(n4528), .Y(n4476) );
  CLKBUFX3 U592 ( .A(n4528), .Y(n4475) );
  CLKBUFX3 U593 ( .A(n4528), .Y(n4474) );
  CLKBUFX3 U594 ( .A(n4529), .Y(n4473) );
  CLKBUFX3 U595 ( .A(n4529), .Y(n4472) );
  CLKBUFX3 U596 ( .A(n4529), .Y(n4471) );
  CLKBUFX3 U597 ( .A(n4529), .Y(n4470) );
  CLKBUFX3 U598 ( .A(n4530), .Y(n4469) );
  CLKBUFX3 U599 ( .A(n4530), .Y(n4468) );
  CLKBUFX3 U600 ( .A(n4530), .Y(n4467) );
  CLKBUFX3 U601 ( .A(n4530), .Y(n4466) );
  CLKBUFX3 U602 ( .A(n4531), .Y(n4465) );
  CLKBUFX3 U603 ( .A(n4531), .Y(n4464) );
  CLKBUFX3 U604 ( .A(n4531), .Y(n4463) );
  CLKBUFX3 U605 ( .A(n4532), .Y(n4461) );
  CLKBUFX3 U606 ( .A(n4532), .Y(n4460) );
  CLKBUFX3 U607 ( .A(n4532), .Y(n4459) );
  CLKBUFX3 U608 ( .A(n4532), .Y(n4458) );
  CLKBUFX3 U609 ( .A(n4533), .Y(n4457) );
  CLKBUFX3 U610 ( .A(n4533), .Y(n4456) );
  CLKBUFX3 U611 ( .A(n4533), .Y(n4455) );
  CLKBUFX3 U612 ( .A(n4533), .Y(n4454) );
  CLKBUFX3 U613 ( .A(n4534), .Y(n4453) );
  CLKBUFX3 U614 ( .A(n4534), .Y(n4452) );
  CLKBUFX3 U615 ( .A(n4534), .Y(n4451) );
  CLKBUFX3 U616 ( .A(n4534), .Y(n4450) );
  INVX3 U617 ( .A(n4444), .Y(n4437) );
  INVX4 U618 ( .A(n4443), .Y(n4438) );
  INVX4 U619 ( .A(n4443), .Y(n4439) );
  CLKBUFX3 U620 ( .A(n4963), .Y(n4406) );
  CLKBUFX3 U621 ( .A(n4963), .Y(n4407) );
  CLKBUFX3 U622 ( .A(n4972), .Y(n4415) );
  CLKBUFX3 U623 ( .A(n4972), .Y(n4416) );
  CLKBUFX3 U624 ( .A(n4967), .Y(n4411) );
  CLKBUFX3 U625 ( .A(n4959), .Y(n4402) );
  CLKBUFX3 U626 ( .A(n4965), .Y(n4408) );
  CLKBUFX3 U627 ( .A(n4958), .Y(n4400) );
  CLKBUFX3 U628 ( .A(n4965), .Y(n4409) );
  CLKBUFX3 U629 ( .A(n4958), .Y(n4401) );
  CLKBUFX3 U630 ( .A(n4969), .Y(n4413) );
  CLKBUFX3 U631 ( .A(n4422), .Y(n4281) );
  CLKBUFX3 U632 ( .A(n4429), .Y(n3757) );
  CLKBUFX3 U633 ( .A(n4429), .Y(n3756) );
  CLKBUFX3 U634 ( .A(n4426), .Y(n4258) );
  CLKBUFX3 U635 ( .A(n4433), .Y(n3733) );
  CLKBUFX3 U636 ( .A(N26), .Y(n4257) );
  CLKBUFX3 U637 ( .A(N21), .Y(n3732) );
  INVX3 U638 ( .A(n4444), .Y(n4436) );
  CLKBUFX3 U639 ( .A(n4518), .Y(n4517) );
  CLKBUFX3 U640 ( .A(n4518), .Y(n4516) );
  CLKBUFX3 U641 ( .A(n4518), .Y(n4515) );
  CLKBUFX3 U642 ( .A(n4518), .Y(n4514) );
  CLKBUFX3 U643 ( .A(n4537), .Y(n4519) );
  CLKBUFX3 U644 ( .A(n4537), .Y(n4520) );
  CLKBUFX3 U645 ( .A(n4536), .Y(n4521) );
  CLKBUFX3 U646 ( .A(n4536), .Y(n4522) );
  CLKBUFX3 U647 ( .A(n4535), .Y(n4523) );
  CLKBUFX3 U648 ( .A(n4535), .Y(n4524) );
  CLKBUFX3 U649 ( .A(n4540), .Y(n4525) );
  CLKBUFX3 U650 ( .A(n4535), .Y(n4526) );
  CLKBUFX3 U651 ( .A(n4540), .Y(n4527) );
  CLKBUFX3 U652 ( .A(n4538), .Y(n4528) );
  CLKBUFX3 U653 ( .A(n4541), .Y(n4529) );
  CLKBUFX3 U654 ( .A(n4536), .Y(n4530) );
  CLKBUFX3 U655 ( .A(n4541), .Y(n4531) );
  CLKBUFX3 U656 ( .A(n4537), .Y(n4532) );
  CLKBUFX3 U657 ( .A(n4538), .Y(n4533) );
  CLKBUFX3 U658 ( .A(n4541), .Y(n4534) );
  CLKBUFX3 U660 ( .A(n4644), .Y(n4367) );
  CLKBUFX3 U661 ( .A(n4644), .Y(n4368) );
  CLKBUFX3 U662 ( .A(n105), .Y(n4307) );
  CLKBUFX3 U663 ( .A(n105), .Y(n4308) );
  CLKBUFX3 U664 ( .A(n106), .Y(n4315) );
  CLKBUFX3 U665 ( .A(n106), .Y(n4316) );
  CLKBUFX3 U666 ( .A(n108), .Y(n4323) );
  CLKBUFX3 U667 ( .A(n108), .Y(n4324) );
  CLKBUFX3 U668 ( .A(n109), .Y(n4331) );
  CLKBUFX3 U669 ( .A(n109), .Y(n4332) );
  CLKBUFX3 U670 ( .A(n110), .Y(n4339) );
  CLKBUFX3 U671 ( .A(n110), .Y(n4340) );
  CLKBUFX3 U672 ( .A(n111), .Y(n4347) );
  CLKBUFX3 U673 ( .A(n111), .Y(n4348) );
  CLKBUFX3 U674 ( .A(n112), .Y(n4355) );
  CLKBUFX3 U675 ( .A(n112), .Y(n4356) );
  NAND2X1 U676 ( .A(n4649), .B(n4650), .Y(n4969) );
  NAND2X1 U677 ( .A(n4645), .B(n4646), .Y(n4961) );
  INVX4 U678 ( .A(n4442), .Y(n4440) );
  CLKBUFX3 U679 ( .A(n4446), .Y(n4443) );
  CLKBUFX3 U680 ( .A(n4446), .Y(n4444) );
  INVX3 U681 ( .A(n4442), .Y(n4441) );
  CLKBUFX3 U682 ( .A(n4967), .Y(n4412) );
  CLKBUFX3 U683 ( .A(n4959), .Y(n4403) );
  CLKBUFX3 U684 ( .A(n4444), .Y(n4445) );
  CLKBUFX3 U685 ( .A(n4638), .Y(n4363) );
  NOR4X1 U686 ( .A(N26), .B(n4426), .C(N24), .D(N23), .Y(n187) );
  NOR4X1 U687 ( .A(n4422), .B(N21), .C(n4433), .D(N19), .Y(n186) );
  CLKINVX1 U688 ( .A(ALUOp[2]), .Y(n4988) );
  CLKBUFX3 U689 ( .A(n4539), .Y(n4537) );
  CLKBUFX3 U690 ( .A(n4539), .Y(n4536) );
  CLKBUFX3 U691 ( .A(n4540), .Y(n4535) );
  CLKBUFX3 U692 ( .A(n4538), .Y(n4518) );
  CLKBUFX3 U693 ( .A(n4539), .Y(n4538) );
  CLKINVX1 U694 ( .A(EX_RegWriteData[0]), .Y(n4955) );
  CLKINVX1 U695 ( .A(EX_RegWriteData[29]), .Y(n4682) );
  CLKINVX1 U696 ( .A(EX_RegWriteData[17]), .Y(n4802) );
  CLKINVX1 U697 ( .A(EX_RegWriteData[16]), .Y(n4793) );
  CLKINVX1 U698 ( .A(EX_RegWriteData[18]), .Y(n4775) );
  CLKINVX1 U699 ( .A(EX_RegWriteData[20]), .Y(n4753) );
  CLKINVX1 U700 ( .A(EX_RegWriteData[23]), .Y(n4744) );
  CLKINVX1 U701 ( .A(EX_RegWriteData[25]), .Y(n4722) );
  CLKINVX1 U702 ( .A(EX_RegWriteData[24]), .Y(n4713) );
  CLKINVX1 U703 ( .A(EX_RegWriteData[27]), .Y(n4704) );
  CLKINVX1 U704 ( .A(EX_RegWriteData[1]), .Y(n4971) );
  CLKINVX1 U705 ( .A(EX_RegWriteData[3]), .Y(n4946) );
  CLKINVX1 U706 ( .A(EX_RegWriteData[2]), .Y(n4937) );
  CLKINVX1 U707 ( .A(EX_RegWriteData[5]), .Y(n4925) );
  CLKINVX1 U708 ( .A(EX_RegWriteData[4]), .Y(n4916) );
  CLKINVX1 U709 ( .A(EX_RegWriteData[7]), .Y(n4907) );
  CLKINVX1 U710 ( .A(EX_RegWriteData[6]), .Y(n4898) );
  CLKINVX1 U711 ( .A(EX_RegWriteData[9]), .Y(n4886) );
  CLKINVX1 U712 ( .A(EX_RegWriteData[8]), .Y(n4877) );
  CLKINVX1 U713 ( .A(EX_RegWriteData[11]), .Y(n4868) );
  CLKINVX1 U714 ( .A(EX_RegWriteData[10]), .Y(n4859) );
  CLKINVX1 U715 ( .A(EX_RegWriteData[13]), .Y(n4846) );
  CLKINVX1 U716 ( .A(EX_RegWriteData[12]), .Y(n4837) );
  CLKINVX1 U717 ( .A(EX_RegWriteData[15]), .Y(n4828) );
  CLKINVX1 U718 ( .A(EX_RegWriteData[14]), .Y(n4819) );
  CLKINVX1 U719 ( .A(EX_RegWriteData[21]), .Y(n4762) );
  CLKINVX1 U720 ( .A(EX_RegWriteData[22]), .Y(n4735) );
  CLKINVX1 U721 ( .A(EX_RegWriteData[26]), .Y(n4695) );
  CLKINVX1 U722 ( .A(EX_RegWriteData[28]), .Y(n4673) );
  CLKINVX1 U723 ( .A(EX_RegWriteData[19]), .Y(n4784) );
  AND2X2 U725 ( .A(n54), .B(n4574), .Y(n105) );
  AND2X2 U726 ( .A(n66), .B(n4574), .Y(n106) );
  AND2X2 U727 ( .A(n76), .B(n4574), .Y(n108) );
  AND2X2 U728 ( .A(n86), .B(n4574), .Y(n109) );
  AND2X2 U729 ( .A(n97), .B(n4574), .Y(n110) );
  AND2X2 U730 ( .A(n107), .B(n4574), .Y(n111) );
  AND2X2 U731 ( .A(n117), .B(n4574), .Y(n112) );
  CLKINVX1 U732 ( .A(n132), .Y(n4575) );
  CLKBUFX3 U733 ( .A(n113), .Y(n4303) );
  CLKBUFX3 U734 ( .A(n113), .Y(n4304) );
  CLKBUFX3 U735 ( .A(n115), .Y(n4309) );
  CLKBUFX3 U736 ( .A(n115), .Y(n4310) );
  CLKBUFX3 U737 ( .A(n135), .Y(n4311) );
  CLKBUFX3 U738 ( .A(n135), .Y(n4312) );
  CLKBUFX3 U739 ( .A(n126), .Y(n4313) );
  CLKBUFX3 U740 ( .A(n126), .Y(n4314) );
  CLKBUFX3 U741 ( .A(n116), .Y(n4317) );
  CLKBUFX3 U742 ( .A(n116), .Y(n4318) );
  CLKBUFX3 U743 ( .A(n136), .Y(n4319) );
  CLKBUFX3 U744 ( .A(n136), .Y(n4320) );
  CLKBUFX3 U745 ( .A(n127), .Y(n4321) );
  CLKBUFX3 U746 ( .A(n127), .Y(n4322) );
  CLKBUFX3 U747 ( .A(n118), .Y(n4325) );
  CLKBUFX3 U748 ( .A(n118), .Y(n4326) );
  CLKBUFX3 U749 ( .A(n137), .Y(n4327) );
  CLKBUFX3 U750 ( .A(n137), .Y(n4328) );
  CLKBUFX3 U751 ( .A(n128), .Y(n4329) );
  CLKBUFX3 U752 ( .A(n128), .Y(n4330) );
  CLKBUFX3 U753 ( .A(n119), .Y(n4333) );
  CLKBUFX3 U754 ( .A(n119), .Y(n4334) );
  CLKBUFX3 U755 ( .A(n138), .Y(n4335) );
  CLKBUFX3 U756 ( .A(n138), .Y(n4336) );
  CLKBUFX3 U757 ( .A(n129), .Y(n4337) );
  CLKBUFX3 U758 ( .A(n129), .Y(n4338) );
  CLKBUFX3 U759 ( .A(n120), .Y(n4341) );
  CLKBUFX3 U760 ( .A(n120), .Y(n4342) );
  CLKBUFX3 U761 ( .A(n139), .Y(n4343) );
  CLKBUFX3 U762 ( .A(n139), .Y(n4344) );
  CLKBUFX3 U763 ( .A(n130), .Y(n4345) );
  CLKBUFX3 U764 ( .A(n130), .Y(n4346) );
  CLKBUFX3 U765 ( .A(n121), .Y(n4349) );
  CLKBUFX3 U766 ( .A(n121), .Y(n4350) );
  CLKBUFX3 U767 ( .A(n140), .Y(n4351) );
  CLKBUFX3 U768 ( .A(n140), .Y(n4352) );
  CLKBUFX3 U769 ( .A(n131), .Y(n4353) );
  CLKBUFX3 U770 ( .A(n131), .Y(n4354) );
  CLKBUFX3 U771 ( .A(n122), .Y(n4357) );
  CLKBUFX3 U772 ( .A(n122), .Y(n4358) );
  CLKBUFX3 U773 ( .A(n123), .Y(n4359) );
  CLKBUFX3 U774 ( .A(n123), .Y(n4360) );
  CLKBUFX3 U775 ( .A(n125), .Y(n4361) );
  CLKBUFX3 U776 ( .A(n125), .Y(n4362) );
  CLKBUFX3 U777 ( .A(n4952), .Y(n4399) );
  CLKBUFX3 U778 ( .A(n4966), .Y(n4410) );
  CLKBUFX3 U779 ( .A(n4934), .Y(n4397) );
  CLKBUFX3 U780 ( .A(n4943), .Y(n4398) );
  CLKBUFX3 U781 ( .A(n4913), .Y(n4395) );
  CLKBUFX3 U782 ( .A(n4922), .Y(n4396) );
  CLKBUFX3 U783 ( .A(n4895), .Y(n4393) );
  CLKBUFX3 U784 ( .A(n4904), .Y(n4394) );
  CLKBUFX3 U785 ( .A(n4874), .Y(n4391) );
  CLKBUFX3 U786 ( .A(n4883), .Y(n4392) );
  CLKBUFX3 U787 ( .A(n4856), .Y(n4389) );
  CLKBUFX3 U788 ( .A(n4865), .Y(n4390) );
  CLKBUFX3 U789 ( .A(n4834), .Y(n4387) );
  CLKBUFX3 U790 ( .A(n4843), .Y(n4388) );
  CLKBUFX3 U791 ( .A(n4816), .Y(n4385) );
  CLKBUFX3 U792 ( .A(n4825), .Y(n4386) );
  CLKBUFX3 U793 ( .A(n4790), .Y(n4383) );
  CLKBUFX3 U794 ( .A(n4799), .Y(n4384) );
  CLKBUFX3 U795 ( .A(n4772), .Y(n4381) );
  CLKBUFX3 U796 ( .A(n4781), .Y(n4382) );
  CLKBUFX3 U797 ( .A(n4750), .Y(n4379) );
  CLKBUFX3 U798 ( .A(n4759), .Y(n4380) );
  CLKBUFX3 U799 ( .A(n4732), .Y(n4377) );
  CLKBUFX3 U800 ( .A(n4741), .Y(n4378) );
  CLKBUFX3 U801 ( .A(n4710), .Y(n4375) );
  CLKBUFX3 U802 ( .A(n4719), .Y(n4376) );
  CLKBUFX3 U803 ( .A(n4692), .Y(n4373) );
  CLKBUFX3 U804 ( .A(n4701), .Y(n4374) );
  CLKBUFX3 U805 ( .A(n4670), .Y(n4371) );
  CLKBUFX3 U806 ( .A(n4679), .Y(n4372) );
  CLKBUFX3 U807 ( .A(n4652), .Y(n4369) );
  CLKBUFX3 U808 ( .A(n4661), .Y(n4370) );
  CLKBUFX3 U809 ( .A(n114), .Y(n4305) );
  CLKBUFX3 U810 ( .A(n114), .Y(n4306) );
  NAND2X1 U811 ( .A(BrForwardB[1]), .B(n4650), .Y(n4965) );
  NAND2X1 U812 ( .A(BrForwardA[1]), .B(n4646), .Y(n4958) );
  NAND2X1 U813 ( .A(BrForwardB[1]), .B(BrForwardB[0]), .Y(n4967) );
  NAND2X1 U814 ( .A(BrForwardA[1]), .B(BrForwardA[0]), .Y(n4959) );
  NAND2X1 U815 ( .A(BrForwardB[0]), .B(n4649), .Y(n4972) );
  NAND2X1 U816 ( .A(BrForwardA[0]), .B(n4645), .Y(n4963) );
  CLKINVX1 U817 ( .A(BrForwardB[0]), .Y(n4650) );
  CLKINVX1 U818 ( .A(BrForwardA[0]), .Y(n4646) );
  CLKINVX1 U819 ( .A(BrForwardB[1]), .Y(n4649) );
  CLKINVX1 U820 ( .A(BrForwardA[1]), .Y(n4645) );
  CLKBUFX3 U821 ( .A(n4447), .Y(n4442) );
  CLKBUFX3 U822 ( .A(n4448), .Y(n4447) );
  CLKBUFX3 U823 ( .A(n4448), .Y(n4446) );
  CLKINVX1 U824 ( .A(n4430), .Y(n4429) );
  CLKINVX1 U825 ( .A(n4427), .Y(n4426) );
  CLKINVX1 U826 ( .A(n4434), .Y(n4433) );
  CLKINVX1 U827 ( .A(Branch), .Y(n4987) );
  CLKBUFX3 U828 ( .A(n4640), .Y(n4364) );
  CLKBUFX3 U829 ( .A(n4449), .Y(n4539) );
  CLKBUFX3 U830 ( .A(n4449), .Y(n4540) );
  CLKBUFX3 U831 ( .A(n4449), .Y(n4541) );
  OA22X1 U832 ( .A0(n4411), .A1(n4790), .B0(n4409), .B1(n4789), .Y(n4791) );
  CLKINVX1 U833 ( .A(next_RData2[16]), .Y(n4792) );
  OA22X1 U834 ( .A0(n4411), .A1(n4781), .B0(n4409), .B1(n4780), .Y(n4782) );
  CLKINVX1 U835 ( .A(next_RData2[19]), .Y(n4783) );
  OA22X1 U836 ( .A0(n4411), .A1(n4772), .B0(n4409), .B1(n4771), .Y(n4773) );
  CLKINVX1 U837 ( .A(next_RData2[18]), .Y(n4774) );
  OA22X1 U838 ( .A0(n4411), .A1(n4750), .B0(n4408), .B1(n4749), .Y(n4751) );
  OA22X1 U839 ( .A0(n4411), .A1(n4741), .B0(n4408), .B1(n4740), .Y(n4742) );
  CLKINVX1 U840 ( .A(next_RData2[23]), .Y(n4743) );
  OA22X1 U841 ( .A0(n4411), .A1(n4732), .B0(n4408), .B1(n4731), .Y(n4733) );
  CLKINVX1 U842 ( .A(next_RData2[22]), .Y(n4734) );
  OA22X1 U843 ( .A0(n4411), .A1(n4710), .B0(n4408), .B1(n4709), .Y(n4711) );
  CLKINVX1 U844 ( .A(next_RData2[24]), .Y(n4712) );
  OA22X1 U845 ( .A0(n4411), .A1(n4701), .B0(n4408), .B1(n4700), .Y(n4702) );
  CLKINVX1 U846 ( .A(next_RData2[27]), .Y(n4703) );
  OA22X1 U847 ( .A0(n4411), .A1(n4692), .B0(n4408), .B1(n4691), .Y(n4693) );
  CLKINVX1 U848 ( .A(next_RData2[26]), .Y(n4694) );
  OA22X1 U849 ( .A0(n4411), .A1(n4670), .B0(n4408), .B1(n4669), .Y(n4671) );
  CLKINVX1 U850 ( .A(next_RData2[28]), .Y(n4672) );
  OA22X1 U851 ( .A0(n4411), .A1(n4661), .B0(n4408), .B1(n4660), .Y(n4662) );
  CLKINVX1 U852 ( .A(next_RData2[31]), .Y(n4663) );
  OA22X1 U853 ( .A0(n4411), .A1(n4652), .B0(n4408), .B1(n4651), .Y(n4653) );
  CLKINVX1 U854 ( .A(next_RData2[30]), .Y(n4654) );
  OA22X1 U855 ( .A0(n4412), .A1(n4952), .B0(n4408), .B1(n4951), .Y(n4953) );
  OA22X1 U856 ( .A0(n4412), .A1(n4943), .B0(n4965), .B1(n4942), .Y(n4944) );
  CLKINVX1 U857 ( .A(next_RData2[3]), .Y(n4945) );
  OA22X1 U858 ( .A0(n4412), .A1(n4934), .B0(n4409), .B1(n4933), .Y(n4935) );
  OA22X1 U859 ( .A0(n4412), .A1(n4913), .B0(n4965), .B1(n4912), .Y(n4914) );
  CLKINVX1 U860 ( .A(next_RData2[4]), .Y(n4915) );
  OA22X1 U861 ( .A0(n4412), .A1(n4904), .B0(n4965), .B1(n4903), .Y(n4905) );
  CLKINVX1 U862 ( .A(next_RData2[7]), .Y(n4906) );
  OA22X1 U863 ( .A0(n4412), .A1(n4895), .B0(n4409), .B1(n4894), .Y(n4896) );
  CLKINVX1 U864 ( .A(next_RData2[6]), .Y(n4897) );
  OA22X1 U865 ( .A0(n4967), .A1(n4874), .B0(n4409), .B1(n4873), .Y(n4875) );
  CLKINVX1 U866 ( .A(next_RData2[8]), .Y(n4876) );
  OA22X1 U867 ( .A0(n4967), .A1(n4865), .B0(n4409), .B1(n4864), .Y(n4866) );
  CLKINVX1 U868 ( .A(next_RData2[11]), .Y(n4867) );
  OA22X1 U869 ( .A0(n4411), .A1(n4856), .B0(n4409), .B1(n4855), .Y(n4857) );
  CLKINVX1 U870 ( .A(next_RData2[10]), .Y(n4858) );
  OA22X1 U871 ( .A0(n4967), .A1(n4834), .B0(n4409), .B1(n4833), .Y(n4835) );
  CLKINVX1 U872 ( .A(next_RData2[12]), .Y(n4836) );
  OA22X1 U873 ( .A0(n4967), .A1(n4825), .B0(n4409), .B1(n4824), .Y(n4826) );
  CLKINVX1 U874 ( .A(next_RData2[15]), .Y(n4827) );
  OA22X1 U875 ( .A0(n4411), .A1(n4816), .B0(n4409), .B1(n4815), .Y(n4817) );
  CLKINVX1 U876 ( .A(next_RData2[14]), .Y(n4818) );
  OA22X1 U877 ( .A0(n4402), .A1(n4790), .B0(n4401), .B1(n4789), .Y(n4787) );
  CLKINVX1 U878 ( .A(next_RData1[16]), .Y(n4788) );
  OA22X1 U880 ( .A0(n4402), .A1(n4772), .B0(n4401), .B1(n4771), .Y(n4769) );
  CLKINVX1 U881 ( .A(next_RData1[18]), .Y(n4770) );
  OA22X1 U882 ( .A0(n4402), .A1(n4750), .B0(n4401), .B1(n4749), .Y(n4747) );
  OA22X1 U888 ( .A0(n4403), .A1(n4710), .B0(n4400), .B1(n4709), .Y(n4707) );
  CLKINVX1 U889 ( .A(next_RData1[24]), .Y(n4708) );
  OA22X1 U890 ( .A0(n4403), .A1(n4701), .B0(n4401), .B1(n4700), .Y(n4698) );
  CLKINVX1 U891 ( .A(next_RData1[27]), .Y(n4699) );
  OA22X1 U892 ( .A0(n4403), .A1(n4692), .B0(n4958), .B1(n4691), .Y(n4689) );
  CLKINVX1 U893 ( .A(next_RData1[26]), .Y(n4690) );
  OA22X1 U896 ( .A0(n4403), .A1(n4661), .B0(n4958), .B1(n4660), .Y(n4658) );
  CLKINVX1 U897 ( .A(next_RData1[31]), .Y(n4659) );
  OA22X1 U898 ( .A0(n4402), .A1(n4652), .B0(n4400), .B1(n4651), .Y(n4647) );
  CLKINVX1 U899 ( .A(next_RData1[30]), .Y(n4648) );
  OA22X1 U900 ( .A0(n4402), .A1(n4952), .B0(n4400), .B1(n4951), .Y(n4949) );
  CLKINVX1 U901 ( .A(next_RData1[0]), .Y(n4950) );
  OA22X1 U902 ( .A0(n4402), .A1(n4943), .B0(n4400), .B1(n4942), .Y(n4940) );
  OA22X1 U903 ( .A0(n4402), .A1(n4934), .B0(n4400), .B1(n4933), .Y(n4931) );
  OA22X1 U904 ( .A0(n4402), .A1(n4913), .B0(n4400), .B1(n4912), .Y(n4910) );
  OA22X1 U905 ( .A0(n4402), .A1(n4904), .B0(n4400), .B1(n4903), .Y(n4901) );
  OA22X1 U907 ( .A0(n4402), .A1(n4895), .B0(n4400), .B1(n4894), .Y(n4892) );
  CLKINVX1 U908 ( .A(next_RData1[6]), .Y(n4893) );
  OA22X1 U909 ( .A0(n4402), .A1(n4874), .B0(n4400), .B1(n4873), .Y(n4871) );
  CLKINVX1 U910 ( .A(next_RData1[8]), .Y(n4872) );
  OA22X1 U911 ( .A0(n4402), .A1(n4865), .B0(n4400), .B1(n4864), .Y(n4862) );
  CLKINVX1 U912 ( .A(next_RData1[11]), .Y(n4863) );
  OA22X1 U913 ( .A0(n4402), .A1(n4856), .B0(n4400), .B1(n4855), .Y(n4853) );
  CLKINVX1 U914 ( .A(next_RData1[10]), .Y(n4854) );
  OA22X1 U915 ( .A0(n4959), .A1(n4834), .B0(n4401), .B1(n4833), .Y(n4831) );
  OA22X1 U917 ( .A0(n4959), .A1(n4825), .B0(n4401), .B1(n4824), .Y(n4822) );
  OA22X1 U918 ( .A0(n4959), .A1(n4816), .B0(n4401), .B1(n4815), .Y(n4813) );
  OA22X1 U921 ( .A0(n4402), .A1(n4759), .B0(n4401), .B1(n4758), .Y(n4756) );
  OA22X1 U922 ( .A0(n4402), .A1(n4719), .B0(n4401), .B1(n4718), .Y(n4716) );
  OA22X1 U923 ( .A0(n4403), .A1(n4679), .B0(n4400), .B1(n4678), .Y(n4676) );
  XNOR2X1 U924 ( .A(n4974), .B(n4973), .Y(n4975) );
  OA22X1 U925 ( .A0(n4959), .A1(n4966), .B0(n4401), .B1(n4964), .Y(n4960) );
  OA22X1 U926 ( .A0(n4402), .A1(n4922), .B0(n4400), .B1(n4921), .Y(n4919) );
  OA22X1 U927 ( .A0(n4402), .A1(n4883), .B0(n4400), .B1(n4882), .Y(n4880) );
  OA22X1 U928 ( .A0(n4959), .A1(n4843), .B0(n4401), .B1(n4842), .Y(n4840) );
  CLKINVX1 U932 ( .A(next_RData1[5]), .Y(n4920) );
  CLKINVX1 U933 ( .A(next_RData1[9]), .Y(n4881) );
  CLKINVX1 U934 ( .A(next_RData1[13]), .Y(n4841) );
  CLKINVX1 U935 ( .A(next_RData2[17]), .Y(n4801) );
  CLKINVX1 U936 ( .A(next_RData2[25]), .Y(n4721) );
  CLKINVX1 U937 ( .A(next_RData2[29]), .Y(n4681) );
  CLKINVX1 U938 ( .A(next_RData2[5]), .Y(n4924) );
  CLKINVX1 U939 ( .A(next_RData2[9]), .Y(n4885) );
  CLKINVX1 U940 ( .A(next_RData2[13]), .Y(n4845) );
  NAND3BX1 U941 ( .AN(n4419), .B(n4420), .C(n4983), .Y(n4644) );
  CLKINVX1 U942 ( .A(EX_RegWriteData[31]), .Y(n4664) );
  NAND2X1 U943 ( .A(n104), .B(n93), .Y(n132) );
  CLKBUFX3 U944 ( .A(n191), .Y(n4420) );
  INVX3 U945 ( .A(n4419), .Y(n4417) );
  AND2X2 U947 ( .A(n54), .B(n53), .Y(n113) );
  AND2X2 U948 ( .A(n54), .B(n57), .Y(n114) );
  AND2X2 U949 ( .A(n66), .B(n65), .Y(n115) );
  AND2X2 U950 ( .A(n76), .B(n65), .Y(n116) );
  AND2X2 U951 ( .A(n86), .B(n65), .Y(n118) );
  AND2X2 U952 ( .A(n97), .B(n65), .Y(n119) );
  AND2X2 U953 ( .A(n107), .B(n65), .Y(n120) );
  AND2X2 U954 ( .A(n117), .B(n65), .Y(n121) );
  AND2X2 U955 ( .A(n65), .B(n4575), .Y(n122) );
  AND2X2 U956 ( .A(n53), .B(n4575), .Y(n123) );
  AND2X2 U957 ( .A(n57), .B(n4575), .Y(n125) );
  AND2X2 U958 ( .A(n66), .B(n57), .Y(n126) );
  AND2X2 U959 ( .A(n76), .B(n57), .Y(n127) );
  AND2X2 U960 ( .A(n86), .B(n57), .Y(n128) );
  AND2X2 U961 ( .A(n97), .B(n57), .Y(n129) );
  AND2X2 U962 ( .A(n107), .B(n57), .Y(n130) );
  AND2X2 U963 ( .A(n117), .B(n57), .Y(n131) );
  AND2X2 U964 ( .A(n66), .B(n53), .Y(n135) );
  AND2X2 U965 ( .A(n76), .B(n53), .Y(n136) );
  AND2X2 U966 ( .A(n86), .B(n53), .Y(n137) );
  AND2X2 U967 ( .A(n97), .B(n53), .Y(n138) );
  AND2X2 U968 ( .A(n107), .B(n53), .Y(n139) );
  AND2X2 U969 ( .A(n117), .B(n53), .Y(n140) );
  AND2X2 U970 ( .A(n104), .B(n83), .Y(n117) );
  AND2X2 U971 ( .A(n73), .B(n61), .Y(n66) );
  AND2X2 U972 ( .A(n83), .B(n61), .Y(n76) );
  AND2X2 U973 ( .A(n93), .B(n61), .Y(n86) );
  AND2X2 U974 ( .A(n104), .B(n62), .Y(n97) );
  AND2X2 U975 ( .A(n104), .B(n73), .Y(n107) );
  AND2X2 U976 ( .A(n61), .B(n62), .Y(n54) );
  CLKBUFX3 U977 ( .A(n191), .Y(n4421) );
  INVX3 U978 ( .A(n4419), .Y(n4418) );
  OA22X1 U979 ( .A0(n4412), .A1(n4799), .B0(n4409), .B1(n4798), .Y(n4800) );
  OA22X1 U980 ( .A0(n4411), .A1(n4759), .B0(n4408), .B1(n4758), .Y(n4760) );
  OA22X1 U981 ( .A0(n4411), .A1(n4719), .B0(n4408), .B1(n4718), .Y(n4720) );
  OA22X1 U982 ( .A0(n4411), .A1(n4679), .B0(n4408), .B1(n4678), .Y(n4680) );
  OA22X1 U983 ( .A0(n4412), .A1(n4966), .B0(n4408), .B1(n4964), .Y(n4968) );
  OA22X1 U984 ( .A0(n4412), .A1(n4922), .B0(n4409), .B1(n4921), .Y(n4923) );
  OA22X1 U985 ( .A0(n4411), .A1(n4883), .B0(n4409), .B1(n4882), .Y(n4884) );
  OA22X1 U986 ( .A0(n4967), .A1(n4843), .B0(n4409), .B1(n4842), .Y(n4844) );
  INVX3 U987 ( .A(n172), .Y(n4985) );
  NOR2X1 U988 ( .A(n4436), .B(Bubble), .Y(n181) );
  OR2X1 U989 ( .A(n167), .B(n4437), .Y(n134) );
  CLKINVX1 U990 ( .A(ALUOp[0]), .Y(n4986) );
  CLKBUFX3 U991 ( .A(rst), .Y(n4449) );
  OAI32X4 U992 ( .A0(n4989), .A1(n4987), .A2(equal), .B0(BranchTaken), .B1(
        n4982), .Y(PredictMiss) );
  MX4X1 U993 ( .A(n247), .B(n245), .C(n246), .D(n244), .S0(n3733), .S1(n3738), 
        .Y(n156) );
  MX4X1 U994 ( .A(n263), .B(n261), .C(n262), .D(n260), .S0(n3734), .S1(n3738), 
        .Y(n160) );
  MX4X1 U995 ( .A(n271), .B(n269), .C(n270), .D(n268), .S0(n3734), .S1(n3738), 
        .Y(n162) );
  MX4X1 U996 ( .A(n279), .B(n277), .C(n278), .D(n276), .S0(n3734), .S1(n3738), 
        .Y(n164) );
  MX4X1 U999 ( .A(n295), .B(n293), .C(n294), .D(n292), .S0(n3734), .S1(n3738), 
        .Y(n173) );
  MX4X1 U1000 ( .A(n303), .B(n301), .C(n302), .D(n300), .S0(n3734), .S1(n3738), 
        .Y(n175) );
  MX4X1 U1001 ( .A(n335), .B(n333), .C(n334), .D(n332), .S0(N20), .S1(n3739), 
        .Y(n197) );
  MX4X1 U1002 ( .A(n343), .B(n341), .C(n342), .D(n340), .S0(N20), .S1(n3739), 
        .Y(n199) );
  MX4X1 U1003 ( .A(n359), .B(n357), .C(n358), .D(n356), .S0(n3735), .S1(N19), 
        .Y(n203) );
  MXI2X1 U1004 ( .A(n205), .B(n206), .S0(N21), .Y(N132) );
  MX4X1 U1005 ( .A(n399), .B(n397), .C(n398), .D(n396), .S0(n3735), .S1(N19), 
        .Y(n213) );
  MX4X1 U1006 ( .A(n423), .B(n421), .C(n422), .D(n420), .S0(n3736), .S1(N19), 
        .Y(n219) );
  MX4X1 U1007 ( .A(n375), .B(n373), .C(n374), .D(n372), .S0(n3735), .S1(N19), 
        .Y(n207) );
  MX4X1 U1008 ( .A(n455), .B(n453), .C(n454), .D(n452), .S0(n3737), .S1(n3740), 
        .Y(n228) );
  MX4X1 U1009 ( .A(n487), .B(n485), .C(n486), .D(n484), .S0(n3737), .S1(n3740), 
        .Y(n236) );
  MX4X1 U1010 ( .A(n495), .B(n493), .C(n494), .D(n492), .S0(n3737), .S1(n3740), 
        .Y(n238) );
  MX4X1 U1011 ( .A(n3860), .B(n3858), .C(n3859), .D(n3857), .S0(n4259), .S1(
        n4262), .Y(n3782) );
  MXI4X1 U1012 ( .A(\regfile[16][2] ), .B(\regfile[17][2] ), .C(
        \regfile[18][2] ), .D(\regfile[19][2] ), .S0(n4291), .S1(n4278), .Y(
        n3860) );
  MXI4X1 U1013 ( .A(\regfile[24][2] ), .B(\regfile[25][2] ), .C(
        \regfile[26][2] ), .D(\regfile[27][2] ), .S0(n4291), .S1(n4276), .Y(
        n3858) );
  MXI4X1 U1014 ( .A(\regfile[28][2] ), .B(\regfile[29][2] ), .C(
        \regfile[30][2] ), .D(\regfile[31][2] ), .S0(n4291), .S1(n4279), .Y(
        n3857) );
  MX4X1 U1015 ( .A(n3868), .B(n3866), .C(n3867), .D(n3865), .S0(n4259), .S1(
        n4262), .Y(n3784) );
  MXI4X1 U1016 ( .A(\regfile[16][3] ), .B(\regfile[17][3] ), .C(
        \regfile[18][3] ), .D(\regfile[19][3] ), .S0(n4292), .S1(n4271), .Y(
        n3868) );
  MXI4X1 U1017 ( .A(\regfile[24][3] ), .B(\regfile[25][3] ), .C(
        \regfile[26][3] ), .D(\regfile[27][3] ), .S0(n4291), .S1(n4271), .Y(
        n3866) );
  MXI4X1 U1018 ( .A(\regfile[28][3] ), .B(\regfile[29][3] ), .C(
        \regfile[30][3] ), .D(\regfile[31][3] ), .S0(n4291), .S1(n4271), .Y(
        n3865) );
  MX4X1 U1019 ( .A(n3876), .B(n3874), .C(n3875), .D(n3873), .S0(n4259), .S1(
        n4262), .Y(n3786) );
  MXI4X1 U1020 ( .A(\regfile[16][4] ), .B(\regfile[17][4] ), .C(
        \regfile[18][4] ), .D(\regfile[19][4] ), .S0(n4292), .S1(n4271), .Y(
        n3876) );
  MXI4X1 U1021 ( .A(\regfile[24][4] ), .B(\regfile[25][4] ), .C(
        \regfile[26][4] ), .D(\regfile[27][4] ), .S0(n4292), .S1(n4271), .Y(
        n3874) );
  MXI4X1 U1022 ( .A(\regfile[28][4] ), .B(\regfile[29][4] ), .C(
        \regfile[30][4] ), .D(\regfile[31][4] ), .S0(n4292), .S1(n4271), .Y(
        n3873) );
  MX4X1 U1023 ( .A(n3884), .B(n3882), .C(n3883), .D(n3881), .S0(n4259), .S1(
        n4262), .Y(n3788) );
  MXI4X1 U1024 ( .A(\regfile[16][5] ), .B(\regfile[17][5] ), .C(
        \regfile[18][5] ), .D(\regfile[19][5] ), .S0(n4292), .S1(n4271), .Y(
        n3884) );
  MXI4X1 U1025 ( .A(\regfile[24][5] ), .B(\regfile[25][5] ), .C(
        \regfile[26][5] ), .D(\regfile[27][5] ), .S0(n4292), .S1(n4271), .Y(
        n3882) );
  MXI4X1 U1026 ( .A(\regfile[28][5] ), .B(\regfile[29][5] ), .C(
        \regfile[30][5] ), .D(\regfile[31][5] ), .S0(n4292), .S1(n4271), .Y(
        n3881) );
  MX4X1 U1027 ( .A(n3892), .B(n3890), .C(n3891), .D(n3889), .S0(n4259), .S1(
        n4262), .Y(n3790) );
  MXI4X1 U1028 ( .A(\regfile[16][6] ), .B(\regfile[17][6] ), .C(
        \regfile[18][6] ), .D(\regfile[19][6] ), .S0(n4293), .S1(n4272), .Y(
        n3892) );
  MXI4X1 U1029 ( .A(\regfile[24][6] ), .B(\regfile[25][6] ), .C(
        \regfile[26][6] ), .D(\regfile[27][6] ), .S0(n4293), .S1(n4272), .Y(
        n3890) );
  MXI4X1 U1030 ( .A(\regfile[28][6] ), .B(\regfile[29][6] ), .C(
        \regfile[30][6] ), .D(\regfile[31][6] ), .S0(n4293), .S1(n4271), .Y(
        n3889) );
  MX4X1 U1031 ( .A(n3900), .B(n3898), .C(n3899), .D(n3897), .S0(n4259), .S1(
        n4262), .Y(n3792) );
  MXI4X1 U1032 ( .A(\regfile[16][7] ), .B(\regfile[17][7] ), .C(
        \regfile[18][7] ), .D(\regfile[19][7] ), .S0(n4293), .S1(n4272), .Y(
        n3900) );
  MXI4X1 U1033 ( .A(\regfile[24][7] ), .B(\regfile[25][7] ), .C(
        \regfile[26][7] ), .D(\regfile[27][7] ), .S0(n4293), .S1(n4272), .Y(
        n3898) );
  MXI4X1 U1034 ( .A(\regfile[28][7] ), .B(\regfile[29][7] ), .C(
        \regfile[30][7] ), .D(\regfile[31][7] ), .S0(n4293), .S1(n4272), .Y(
        n3897) );
  MX4X1 U1035 ( .A(n3908), .B(n3906), .C(n3907), .D(n3905), .S0(N25), .S1(N24), 
        .Y(n3794) );
  MXI4X1 U1036 ( .A(\regfile[16][8] ), .B(\regfile[17][8] ), .C(
        \regfile[18][8] ), .D(\regfile[19][8] ), .S0(n4294), .S1(n4272), .Y(
        n3908) );
  MXI4X1 U1037 ( .A(\regfile[24][8] ), .B(\regfile[25][8] ), .C(
        \regfile[26][8] ), .D(\regfile[27][8] ), .S0(n4294), .S1(n4272), .Y(
        n3906) );
  MXI4X1 U1038 ( .A(\regfile[28][8] ), .B(\regfile[29][8] ), .C(
        \regfile[30][8] ), .D(\regfile[31][8] ), .S0(n4297), .S1(n4275), .Y(
        n3905) );
  MX4X1 U1039 ( .A(n3916), .B(n3914), .C(n3915), .D(n3913), .S0(N25), .S1(
        n4264), .Y(n3796) );
  MXI4X1 U1040 ( .A(\regfile[16][9] ), .B(\regfile[17][9] ), .C(
        \regfile[18][9] ), .D(\regfile[19][9] ), .S0(n4294), .S1(n4273), .Y(
        n3916) );
  MXI4X1 U1041 ( .A(\regfile[24][9] ), .B(\regfile[25][9] ), .C(
        \regfile[26][9] ), .D(\regfile[27][9] ), .S0(n4294), .S1(n4273), .Y(
        n3914) );
  MXI4X1 U1042 ( .A(\regfile[28][9] ), .B(\regfile[29][9] ), .C(
        \regfile[30][9] ), .D(\regfile[31][9] ), .S0(n4294), .S1(n4272), .Y(
        n3913) );
  MXI4X1 U1044 ( .A(\regfile[16][10] ), .B(\regfile[17][10] ), .C(
        \regfile[18][10] ), .D(\regfile[19][10] ), .S0(n4295), .S1(n4273), .Y(
        n3924) );
  MXI4X1 U1045 ( .A(\regfile[24][10] ), .B(\regfile[25][10] ), .C(
        \regfile[26][10] ), .D(\regfile[27][10] ), .S0(n4295), .S1(n4273), .Y(
        n3922) );
  MXI4X1 U1046 ( .A(\regfile[28][10] ), .B(\regfile[29][10] ), .C(
        \regfile[30][10] ), .D(\regfile[31][10] ), .S0(n4295), .S1(n4273), .Y(
        n3921) );
  MX4X1 U1047 ( .A(n3932), .B(n3930), .C(n3931), .D(n3929), .S0(N25), .S1(N24), 
        .Y(n3800) );
  MXI4X1 U1048 ( .A(\regfile[16][11] ), .B(\regfile[17][11] ), .C(
        \regfile[18][11] ), .D(\regfile[19][11] ), .S0(n4295), .S1(n4273), .Y(
        n3932) );
  MXI4X1 U1049 ( .A(\regfile[24][11] ), .B(\regfile[25][11] ), .C(
        \regfile[26][11] ), .D(\regfile[27][11] ), .S0(n4295), .S1(n4273), .Y(
        n3930) );
  MXI4X1 U1050 ( .A(\regfile[28][11] ), .B(\regfile[29][11] ), .C(
        \regfile[30][11] ), .D(\regfile[31][11] ), .S0(n4295), .S1(n4273), .Y(
        n3929) );
  MXI4X1 U1052 ( .A(\regfile[16][12] ), .B(\regfile[17][12] ), .C(
        \regfile[18][12] ), .D(\regfile[19][12] ), .S0(n4296), .S1(n4266), .Y(
        n3940) );
  MXI4X1 U1053 ( .A(\regfile[24][12] ), .B(\regfile[25][12] ), .C(
        \regfile[26][12] ), .D(\regfile[27][12] ), .S0(n4296), .S1(n4273), .Y(
        n3938) );
  MXI4X1 U1054 ( .A(\regfile[28][12] ), .B(\regfile[29][12] ), .C(
        \regfile[30][12] ), .D(\regfile[31][12] ), .S0(n4296), .S1(n4273), .Y(
        n3937) );
  MX4X1 U1055 ( .A(n3948), .B(n3946), .C(n3947), .D(n3945), .S0(N25), .S1(N24), 
        .Y(n3804) );
  MXI4X1 U1056 ( .A(\regfile[16][13] ), .B(\regfile[17][13] ), .C(
        \regfile[18][13] ), .D(\regfile[19][13] ), .S0(n4296), .S1(n4272), .Y(
        n3948) );
  MXI4X1 U1057 ( .A(\regfile[24][13] ), .B(\regfile[25][13] ), .C(
        \regfile[26][13] ), .D(\regfile[27][13] ), .S0(n4296), .S1(n4276), .Y(
        n3946) );
  MXI4X1 U1058 ( .A(\regfile[28][13] ), .B(\regfile[29][13] ), .C(
        \regfile[30][13] ), .D(\regfile[31][13] ), .S0(n4296), .S1(n4274), .Y(
        n3945) );
  MX4X1 U1059 ( .A(n3956), .B(n3954), .C(n3955), .D(n3953), .S0(N25), .S1(
        n4263), .Y(n3806) );
  MXI4X1 U1060 ( .A(\regfile[16][14] ), .B(\regfile[17][14] ), .C(
        \regfile[18][14] ), .D(\regfile[19][14] ), .S0(n4297), .S1(n4268), .Y(
        n3956) );
  MXI4X1 U1061 ( .A(\regfile[24][14] ), .B(\regfile[25][14] ), .C(
        \regfile[26][14] ), .D(\regfile[27][14] ), .S0(n4297), .S1(n4267), .Y(
        n3954) );
  MXI4X1 U1062 ( .A(\regfile[28][14] ), .B(\regfile[29][14] ), .C(
        \regfile[30][14] ), .D(\regfile[31][14] ), .S0(n4296), .S1(n4280), .Y(
        n3953) );
  MX4X1 U1063 ( .A(n3964), .B(n3962), .C(n3963), .D(n3961), .S0(N25), .S1(
        n4263), .Y(n3808) );
  MXI4X1 U1064 ( .A(\regfile[16][15] ), .B(\regfile[17][15] ), .C(
        \regfile[18][15] ), .D(\regfile[19][15] ), .S0(n4297), .S1(n4273), .Y(
        n3964) );
  MXI4X1 U1065 ( .A(\regfile[24][15] ), .B(\regfile[25][15] ), .C(
        \regfile[26][15] ), .D(\regfile[27][15] ), .S0(n4297), .S1(n4272), .Y(
        n3962) );
  MXI4X1 U1066 ( .A(\regfile[28][15] ), .B(\regfile[29][15] ), .C(
        \regfile[30][15] ), .D(\regfile[31][15] ), .S0(n4297), .S1(n4266), .Y(
        n3961) );
  MX4X1 U1067 ( .A(n3972), .B(n3970), .C(n3971), .D(n3969), .S0(N25), .S1(
        n4263), .Y(n3810) );
  MXI4X1 U1068 ( .A(\regfile[16][16] ), .B(\regfile[17][16] ), .C(
        \regfile[18][16] ), .D(\regfile[19][16] ), .S0(n4283), .S1(n4269), .Y(
        n3972) );
  MXI4X1 U1069 ( .A(\regfile[24][16] ), .B(\regfile[25][16] ), .C(
        \regfile[26][16] ), .D(\regfile[27][16] ), .S0(n4283), .S1(n4270), .Y(
        n3970) );
  MXI4X1 U1070 ( .A(\regfile[28][16] ), .B(\regfile[29][16] ), .C(
        \regfile[30][16] ), .D(\regfile[31][16] ), .S0(n4283), .S1(n4275), .Y(
        n3969) );
  MX4X1 U1071 ( .A(n3980), .B(n3978), .C(n3979), .D(n3977), .S0(N25), .S1(
        n4263), .Y(n3812) );
  MXI4X1 U1072 ( .A(\regfile[16][17] ), .B(\regfile[17][17] ), .C(
        \regfile[18][17] ), .D(\regfile[19][17] ), .S0(n4283), .S1(n4280), .Y(
        n3980) );
  MXI4X1 U1073 ( .A(\regfile[24][17] ), .B(\regfile[25][17] ), .C(
        \regfile[26][17] ), .D(\regfile[27][17] ), .S0(n4283), .S1(n4270), .Y(
        n3978) );
  MXI4X1 U1074 ( .A(\regfile[28][17] ), .B(\regfile[29][17] ), .C(
        \regfile[30][17] ), .D(\regfile[31][17] ), .S0(n4283), .S1(n4268), .Y(
        n3977) );
  MX4X1 U1075 ( .A(n3988), .B(n3986), .C(n3987), .D(n3985), .S0(N25), .S1(
        n4263), .Y(n3814) );
  MXI4X1 U1076 ( .A(\regfile[16][18] ), .B(\regfile[17][18] ), .C(
        \regfile[18][18] ), .D(\regfile[19][18] ), .S0(n4284), .S1(n4278), .Y(
        n3988) );
  MXI4X1 U1077 ( .A(\regfile[24][18] ), .B(\regfile[25][18] ), .C(
        \regfile[26][18] ), .D(\regfile[27][18] ), .S0(n4284), .S1(n4279), .Y(
        n3986) );
  MXI4X1 U1078 ( .A(\regfile[28][18] ), .B(\regfile[29][18] ), .C(
        \regfile[30][18] ), .D(\regfile[31][18] ), .S0(n4283), .S1(n4280), .Y(
        n3985) );
  MX4X1 U1079 ( .A(n3996), .B(n3994), .C(n3995), .D(n3993), .S0(N25), .S1(
        n4263), .Y(n3816) );
  MXI4X1 U1080 ( .A(\regfile[16][19] ), .B(\regfile[17][19] ), .C(
        \regfile[18][19] ), .D(\regfile[19][19] ), .S0(n4284), .S1(n4276), .Y(
        n3996) );
  MXI4X1 U1081 ( .A(\regfile[24][19] ), .B(\regfile[25][19] ), .C(
        \regfile[26][19] ), .D(\regfile[27][19] ), .S0(n4284), .S1(n4277), .Y(
        n3994) );
  MXI4X1 U1082 ( .A(\regfile[28][19] ), .B(\regfile[29][19] ), .C(
        \regfile[30][19] ), .D(\regfile[31][19] ), .S0(n4284), .S1(n4275), .Y(
        n3993) );
  MXI4X1 U1084 ( .A(\regfile[16][20] ), .B(\regfile[17][20] ), .C(
        \regfile[18][20] ), .D(\regfile[19][20] ), .S0(n4285), .S1(n4267), .Y(
        n4004) );
  MXI4X1 U1085 ( .A(\regfile[24][20] ), .B(\regfile[25][20] ), .C(
        \regfile[26][20] ), .D(\regfile[27][20] ), .S0(n4284), .S1(n4267), .Y(
        n4002) );
  MXI4X1 U1086 ( .A(\regfile[28][20] ), .B(\regfile[29][20] ), .C(
        \regfile[30][20] ), .D(\regfile[31][20] ), .S0(n4284), .S1(n4267), .Y(
        n4001) );
  MXI4X1 U1088 ( .A(\regfile[16][21] ), .B(\regfile[17][21] ), .C(
        \regfile[18][21] ), .D(\regfile[19][21] ), .S0(n4285), .S1(n4266), .Y(
        n4012) );
  MXI4X1 U1089 ( .A(\regfile[24][21] ), .B(\regfile[25][21] ), .C(
        \regfile[26][21] ), .D(\regfile[27][21] ), .S0(n4285), .S1(n4267), .Y(
        n4010) );
  MXI4X1 U1090 ( .A(\regfile[28][21] ), .B(\regfile[29][21] ), .C(
        \regfile[30][21] ), .D(\regfile[31][21] ), .S0(n4285), .S1(n4266), .Y(
        n4009) );
  MX4X1 U1091 ( .A(n4020), .B(n4018), .C(n4019), .D(n4017), .S0(n4261), .S1(
        n4264), .Y(n3822) );
  MXI4X1 U1092 ( .A(\regfile[16][22] ), .B(\regfile[17][22] ), .C(
        \regfile[18][22] ), .D(\regfile[19][22] ), .S0(n4286), .S1(n4279), .Y(
        n4020) );
  MXI4X1 U1093 ( .A(\regfile[24][22] ), .B(\regfile[25][22] ), .C(
        \regfile[26][22] ), .D(\regfile[27][22] ), .S0(n4285), .S1(n4276), .Y(
        n4018) );
  MXI4X1 U1094 ( .A(\regfile[28][22] ), .B(\regfile[29][22] ), .C(
        \regfile[30][22] ), .D(\regfile[31][22] ), .S0(n4285), .S1(n4276), .Y(
        n4017) );
  MX4X1 U1095 ( .A(n4028), .B(n4026), .C(n4027), .D(n4025), .S0(n4261), .S1(
        n4264), .Y(n3824) );
  MXI4X1 U1096 ( .A(\regfile[16][23] ), .B(\regfile[17][23] ), .C(
        \regfile[18][23] ), .D(\regfile[19][23] ), .S0(n4286), .S1(n4268), .Y(
        n4028) );
  MXI4X1 U1097 ( .A(\regfile[24][23] ), .B(\regfile[25][23] ), .C(
        \regfile[26][23] ), .D(\regfile[27][23] ), .S0(n4286), .S1(n4275), .Y(
        n4026) );
  MXI4X1 U1098 ( .A(\regfile[28][23] ), .B(\regfile[29][23] ), .C(
        \regfile[30][23] ), .D(\regfile[31][23] ), .S0(n4286), .S1(n4276), .Y(
        n4025) );
  MX4X1 U1099 ( .A(n4036), .B(n4034), .C(n4035), .D(n4033), .S0(n4261), .S1(
        n4264), .Y(n3826) );
  MXI4X1 U1100 ( .A(\regfile[16][24] ), .B(\regfile[17][24] ), .C(
        \regfile[18][24] ), .D(\regfile[19][24] ), .S0(n4287), .S1(n4269), .Y(
        n4036) );
  MXI4X1 U1101 ( .A(\regfile[24][24] ), .B(\regfile[25][24] ), .C(
        \regfile[26][24] ), .D(\regfile[27][24] ), .S0(n4286), .S1(n4279), .Y(
        n4034) );
  MXI4X1 U1102 ( .A(\regfile[28][24] ), .B(\regfile[29][24] ), .C(
        \regfile[30][24] ), .D(\regfile[31][24] ), .S0(n4286), .S1(n4280), .Y(
        n4033) );
  MX4X1 U1103 ( .A(n4044), .B(n4042), .C(n4043), .D(n4041), .S0(n4261), .S1(
        n4264), .Y(n3828) );
  MXI4X1 U1104 ( .A(\regfile[16][25] ), .B(\regfile[17][25] ), .C(
        \regfile[18][25] ), .D(\regfile[19][25] ), .S0(n4287), .S1(n4280), .Y(
        n4044) );
  MXI4X1 U1105 ( .A(\regfile[24][25] ), .B(\regfile[25][25] ), .C(
        \regfile[26][25] ), .D(\regfile[27][25] ), .S0(n4287), .S1(n4276), .Y(
        n4042) );
  MXI4X1 U1106 ( .A(\regfile[28][25] ), .B(\regfile[29][25] ), .C(
        \regfile[30][25] ), .D(\regfile[31][25] ), .S0(n4287), .S1(n4275), .Y(
        n4041) );
  MX4X1 U1107 ( .A(n4052), .B(n4050), .C(n4051), .D(n4049), .S0(N25), .S1(
        n4265), .Y(n3830) );
  MXI4X1 U1108 ( .A(\regfile[16][26] ), .B(\regfile[17][26] ), .C(
        \regfile[18][26] ), .D(\regfile[19][26] ), .S0(n4287), .S1(n4267), .Y(
        n4052) );
  MXI4X1 U1109 ( .A(\regfile[24][26] ), .B(\regfile[25][26] ), .C(
        \regfile[26][26] ), .D(\regfile[27][26] ), .S0(n4287), .S1(n4267), .Y(
        n4050) );
  MXI4X1 U1110 ( .A(\regfile[28][26] ), .B(\regfile[29][26] ), .C(
        \regfile[30][26] ), .D(\regfile[31][26] ), .S0(n4287), .S1(n4267), .Y(
        n4049) );
  MX4X1 U1111 ( .A(n4060), .B(n4058), .C(n4059), .D(n4057), .S0(n4258), .S1(
        n4265), .Y(n3832) );
  MXI4X1 U1112 ( .A(\regfile[16][27] ), .B(\regfile[17][27] ), .C(
        \regfile[18][27] ), .D(\regfile[19][27] ), .S0(n4288), .S1(n4267), .Y(
        n4060) );
  MXI4X1 U1113 ( .A(\regfile[24][27] ), .B(\regfile[25][27] ), .C(
        \regfile[26][27] ), .D(\regfile[27][27] ), .S0(n4288), .S1(n4267), .Y(
        n4058) );
  MXI4X1 U1114 ( .A(\regfile[28][27] ), .B(\regfile[29][27] ), .C(
        \regfile[30][27] ), .D(\regfile[31][27] ), .S0(n4288), .S1(n4276), .Y(
        n4057) );
  MX4X1 U1115 ( .A(n4068), .B(n4066), .C(n4067), .D(n4065), .S0(n4426), .S1(
        n4265), .Y(n3834) );
  MXI4X1 U1116 ( .A(\regfile[16][28] ), .B(\regfile[17][28] ), .C(
        \regfile[18][28] ), .D(\regfile[19][28] ), .S0(n4288), .S1(n4280), .Y(
        n4068) );
  MXI4X1 U1117 ( .A(\regfile[24][28] ), .B(\regfile[25][28] ), .C(
        \regfile[26][28] ), .D(\regfile[27][28] ), .S0(n4288), .S1(n4275), .Y(
        n4066) );
  MXI4X1 U1118 ( .A(\regfile[28][28] ), .B(\regfile[29][28] ), .C(
        \regfile[30][28] ), .D(\regfile[31][28] ), .S0(n4288), .S1(n4275), .Y(
        n4065) );
  MX4X1 U1119 ( .A(n4076), .B(n4074), .C(n4075), .D(n4073), .S0(N25), .S1(
        n4265), .Y(n3836) );
  MXI4X1 U1120 ( .A(\regfile[16][29] ), .B(\regfile[17][29] ), .C(
        \regfile[18][29] ), .D(\regfile[19][29] ), .S0(n4289), .S1(n4269), .Y(
        n4076) );
  MXI4X1 U1121 ( .A(\regfile[24][29] ), .B(\regfile[25][29] ), .C(
        \regfile[26][29] ), .D(\regfile[27][29] ), .S0(n4289), .S1(n4274), .Y(
        n4074) );
  MXI4X1 U1122 ( .A(\regfile[28][29] ), .B(\regfile[29][29] ), .C(
        \regfile[30][29] ), .D(\regfile[31][29] ), .S0(n4289), .S1(n4279), .Y(
        n4073) );
  MX4X1 U1123 ( .A(n4084), .B(n4082), .C(n4083), .D(n4081), .S0(N25), .S1(
        n4265), .Y(n3838) );
  MXI4X1 U1124 ( .A(\regfile[16][30] ), .B(\regfile[17][30] ), .C(
        \regfile[18][30] ), .D(\regfile[19][30] ), .S0(n4289), .S1(n4274), .Y(
        n4084) );
  MXI4X1 U1125 ( .A(\regfile[24][30] ), .B(\regfile[25][30] ), .C(
        \regfile[26][30] ), .D(\regfile[27][30] ), .S0(n4289), .S1(n4279), .Y(
        n4082) );
  MXI4X1 U1126 ( .A(\regfile[28][30] ), .B(\regfile[29][30] ), .C(
        \regfile[30][30] ), .D(\regfile[31][30] ), .S0(n4289), .S1(n4276), .Y(
        n4081) );
  MXI4X1 U1128 ( .A(\regfile[16][31] ), .B(\regfile[17][31] ), .C(
        \regfile[18][31] ), .D(\regfile[19][31] ), .S0(n4290), .S1(n4271), .Y(
        n4092) );
  MXI4X1 U1129 ( .A(\regfile[24][31] ), .B(\regfile[25][31] ), .C(
        \regfile[26][31] ), .D(\regfile[27][31] ), .S0(n4290), .S1(n4266), .Y(
        n4090) );
  MXI4X1 U1130 ( .A(\regfile[28][31] ), .B(\regfile[29][31] ), .C(
        \regfile[30][31] ), .D(\regfile[31][31] ), .S0(n4290), .S1(n4266), .Y(
        n4089) );
  MX4X1 U1131 ( .A(n259), .B(n257), .C(n258), .D(n256), .S0(n3734), .S1(n3738), 
        .Y(n161) );
  MXI4X1 U1132 ( .A(\regfile[16][2] ), .B(\regfile[17][2] ), .C(
        \regfile[18][2] ), .D(\regfile[19][2] ), .S0(n3766), .S1(n3745), .Y(
        n259) );
  MXI4X1 U1133 ( .A(\regfile[24][2] ), .B(\regfile[25][2] ), .C(
        \regfile[26][2] ), .D(\regfile[27][2] ), .S0(n3766), .S1(n3745), .Y(
        n257) );
  MXI4X1 U1134 ( .A(\regfile[28][2] ), .B(\regfile[29][2] ), .C(
        \regfile[30][2] ), .D(\regfile[31][2] ), .S0(n3766), .S1(n3745), .Y(
        n256) );
  MX4X1 U1135 ( .A(n267), .B(n265), .C(n266), .D(n264), .S0(n3734), .S1(n3738), 
        .Y(n163) );
  MXI4X1 U1136 ( .A(\regfile[16][3] ), .B(\regfile[17][3] ), .C(
        \regfile[18][3] ), .D(\regfile[19][3] ), .S0(n3767), .S1(n3751), .Y(
        n267) );
  MXI4X1 U1137 ( .A(\regfile[24][3] ), .B(\regfile[25][3] ), .C(
        \regfile[26][3] ), .D(\regfile[27][3] ), .S0(n3766), .S1(n3743), .Y(
        n265) );
  MXI4X1 U1138 ( .A(\regfile[28][3] ), .B(\regfile[29][3] ), .C(
        \regfile[30][3] ), .D(\regfile[31][3] ), .S0(n3766), .S1(n3746), .Y(
        n264) );
  MX4X1 U1139 ( .A(n275), .B(n273), .C(n274), .D(n272), .S0(n3734), .S1(n3738), 
        .Y(n165) );
  MXI4X1 U1140 ( .A(\regfile[16][4] ), .B(\regfile[17][4] ), .C(
        \regfile[18][4] ), .D(\regfile[19][4] ), .S0(n3767), .S1(n3746), .Y(
        n275) );
  MXI4X1 U1141 ( .A(\regfile[24][4] ), .B(\regfile[25][4] ), .C(
        \regfile[26][4] ), .D(\regfile[27][4] ), .S0(n3767), .S1(n3755), .Y(
        n273) );
  MXI4X1 U1142 ( .A(\regfile[28][4] ), .B(\regfile[29][4] ), .C(
        \regfile[30][4] ), .D(\regfile[31][4] ), .S0(n3767), .S1(n3753), .Y(
        n272) );
  MXI4X1 U1144 ( .A(\regfile[16][5] ), .B(\regfile[17][5] ), .C(
        \regfile[18][5] ), .D(\regfile[19][5] ), .S0(n3767), .S1(n3751), .Y(
        n283) );
  MXI4X1 U1145 ( .A(\regfile[24][5] ), .B(\regfile[25][5] ), .C(
        \regfile[26][5] ), .D(\regfile[27][5] ), .S0(n3767), .S1(n3753), .Y(
        n281) );
  MXI4X1 U1146 ( .A(\regfile[28][5] ), .B(\regfile[29][5] ), .C(
        \regfile[30][5] ), .D(\regfile[31][5] ), .S0(n3767), .S1(n3755), .Y(
        n280) );
  MX4X1 U1147 ( .A(n291), .B(n289), .C(n290), .D(n288), .S0(n3734), .S1(n3738), 
        .Y(n174) );
  MXI4X1 U1148 ( .A(\regfile[28][6] ), .B(\regfile[29][6] ), .C(
        \regfile[30][6] ), .D(\regfile[31][6] ), .S0(n3768), .S1(n3755), .Y(
        n288) );
  MX4X1 U1149 ( .A(n299), .B(n297), .C(n298), .D(n296), .S0(n3734), .S1(n3738), 
        .Y(n188) );
  MXI4X1 U1150 ( .A(\regfile[24][7] ), .B(\regfile[25][7] ), .C(
        \regfile[26][7] ), .D(\regfile[27][7] ), .S0(n3768), .S1(n3742), .Y(
        n297) );
  MXI4X1 U1151 ( .A(\regfile[28][7] ), .B(\regfile[29][7] ), .C(
        \regfile[30][7] ), .D(\regfile[31][7] ), .S0(n3768), .S1(n3745), .Y(
        n296) );
  MX4X1 U1152 ( .A(n307), .B(n305), .C(n306), .D(n304), .S0(N20), .S1(n3739), 
        .Y(n190) );
  MXI4X1 U1153 ( .A(\regfile[16][8] ), .B(\regfile[17][8] ), .C(
        \regfile[18][8] ), .D(\regfile[19][8] ), .S0(n3769), .S1(n3754), .Y(
        n307) );
  MXI4X1 U1154 ( .A(\regfile[24][8] ), .B(\regfile[25][8] ), .C(
        \regfile[26][8] ), .D(\regfile[27][8] ), .S0(n3769), .S1(n3755), .Y(
        n305) );
  MXI4X1 U1155 ( .A(\regfile[28][8] ), .B(\regfile[29][8] ), .C(
        \regfile[30][8] ), .D(\regfile[31][8] ), .S0(n3772), .S1(n3749), .Y(
        n304) );
  MX4X1 U1156 ( .A(n315), .B(n313), .C(n314), .D(n312), .S0(N20), .S1(n3739), 
        .Y(n194) );
  MXI4X1 U1157 ( .A(\regfile[16][9] ), .B(\regfile[17][9] ), .C(
        \regfile[18][9] ), .D(\regfile[19][9] ), .S0(n3769), .S1(n3747), .Y(
        n315) );
  MXI4X1 U1158 ( .A(\regfile[24][9] ), .B(\regfile[25][9] ), .C(
        \regfile[26][9] ), .D(\regfile[27][9] ), .S0(n3769), .S1(n3747), .Y(
        n313) );
  MXI4X1 U1159 ( .A(\regfile[28][9] ), .B(\regfile[29][9] ), .C(
        \regfile[30][9] ), .D(\regfile[31][9] ), .S0(n3769), .S1(n3743), .Y(
        n312) );
  MX4X1 U1160 ( .A(n323), .B(n321), .C(n322), .D(n320), .S0(N20), .S1(n3739), 
        .Y(n196) );
  MXI4X1 U1161 ( .A(\regfile[16][10] ), .B(\regfile[17][10] ), .C(
        \regfile[18][10] ), .D(\regfile[19][10] ), .S0(n3770), .S1(n3747), .Y(
        n323) );
  MXI4X1 U1162 ( .A(\regfile[24][10] ), .B(\regfile[25][10] ), .C(
        \regfile[26][10] ), .D(\regfile[27][10] ), .S0(n3770), .S1(n3747), .Y(
        n321) );
  MXI4X1 U1163 ( .A(\regfile[28][10] ), .B(\regfile[29][10] ), .C(
        \regfile[30][10] ), .D(\regfile[31][10] ), .S0(n3770), .S1(n3747), .Y(
        n320) );
  MXI4X1 U1164 ( .A(\regfile[16][11] ), .B(\regfile[17][11] ), .C(
        \regfile[18][11] ), .D(\regfile[19][11] ), .S0(n3770), .S1(n3747), .Y(
        n331) );
  MXI4X1 U1165 ( .A(\regfile[24][11] ), .B(\regfile[25][11] ), .C(
        \regfile[26][11] ), .D(\regfile[27][11] ), .S0(n3770), .S1(n3747), .Y(
        n329) );
  MXI4X1 U1166 ( .A(\regfile[28][11] ), .B(\regfile[29][11] ), .C(
        \regfile[30][11] ), .D(\regfile[31][11] ), .S0(n3770), .S1(n3747), .Y(
        n328) );
  MX4X1 U1167 ( .A(n339), .B(n337), .C(n338), .D(n336), .S0(N20), .S1(n3739), 
        .Y(n200) );
  MXI4X1 U1168 ( .A(\regfile[16][12] ), .B(\regfile[17][12] ), .C(
        \regfile[18][12] ), .D(\regfile[19][12] ), .S0(n3771), .S1(n3743), .Y(
        n339) );
  MXI4X1 U1169 ( .A(\regfile[24][12] ), .B(\regfile[25][12] ), .C(
        \regfile[26][12] ), .D(\regfile[27][12] ), .S0(n3771), .S1(n3747), .Y(
        n337) );
  MXI4X1 U1170 ( .A(\regfile[28][12] ), .B(\regfile[29][12] ), .C(
        \regfile[30][12] ), .D(\regfile[31][12] ), .S0(n3771), .S1(n3747), .Y(
        n336) );
  MX4X1 U1171 ( .A(n347), .B(n345), .C(n346), .D(n344), .S0(N20), .S1(n3739), 
        .Y(n202) );
  MXI4X1 U1172 ( .A(\regfile[16][13] ), .B(\regfile[17][13] ), .C(
        \regfile[18][13] ), .D(\regfile[19][13] ), .S0(n3771), .S1(n3743), .Y(
        n347) );
  MXI4X1 U1173 ( .A(\regfile[24][13] ), .B(\regfile[25][13] ), .C(
        \regfile[26][13] ), .D(\regfile[27][13] ), .S0(n3771), .S1(n3752), .Y(
        n345) );
  MXI4X1 U1174 ( .A(\regfile[28][13] ), .B(\regfile[29][13] ), .C(
        \regfile[30][13] ), .D(\regfile[31][13] ), .S0(n3771), .S1(n3753), .Y(
        n344) );
  MX4X1 U1175 ( .A(n355), .B(n353), .C(n354), .D(n352), .S0(n3735), .S1(N19), 
        .Y(n204) );
  MXI4X1 U1176 ( .A(\regfile[16][14] ), .B(\regfile[17][14] ), .C(
        \regfile[18][14] ), .D(\regfile[19][14] ), .S0(n3772), .S1(n3753), .Y(
        n355) );
  MXI4X1 U1177 ( .A(\regfile[24][14] ), .B(\regfile[25][14] ), .C(
        \regfile[26][14] ), .D(\regfile[27][14] ), .S0(n3772), .S1(n3752), .Y(
        n353) );
  MXI4X1 U1178 ( .A(\regfile[28][14] ), .B(\regfile[29][14] ), .C(
        \regfile[30][14] ), .D(\regfile[31][14] ), .S0(n3771), .S1(n3748), .Y(
        n352) );
  MX4X1 U1179 ( .A(n363), .B(n361), .C(n362), .D(n360), .S0(n3735), .S1(n3738), 
        .Y(n206) );
  MXI4X1 U1180 ( .A(\regfile[16][15] ), .B(\regfile[17][15] ), .C(
        \regfile[18][15] ), .D(\regfile[19][15] ), .S0(n3772), .S1(n3755), .Y(
        n363) );
  MXI4X1 U1181 ( .A(\regfile[24][15] ), .B(\regfile[25][15] ), .C(
        \regfile[26][15] ), .D(\regfile[27][15] ), .S0(n3772), .S1(n3754), .Y(
        n361) );
  MXI4X1 U1182 ( .A(\regfile[28][15] ), .B(\regfile[29][15] ), .C(
        \regfile[30][15] ), .D(\regfile[31][15] ), .S0(n3772), .S1(n3751), .Y(
        n360) );
  MX4X1 U1183 ( .A(n371), .B(n369), .C(n370), .D(n368), .S0(n3735), .S1(n3738), 
        .Y(n208) );
  MXI4X1 U1184 ( .A(\regfile[16][16] ), .B(\regfile[17][16] ), .C(
        \regfile[18][16] ), .D(\regfile[19][16] ), .S0(n3758), .S1(n3742), .Y(
        n371) );
  MXI4X1 U1185 ( .A(\regfile[24][16] ), .B(\regfile[25][16] ), .C(
        \regfile[26][16] ), .D(\regfile[27][16] ), .S0(n3758), .S1(n3743), .Y(
        n369) );
  MXI4X1 U1186 ( .A(\regfile[28][16] ), .B(\regfile[29][16] ), .C(
        \regfile[30][16] ), .D(\regfile[31][16] ), .S0(n3758), .S1(n3755), .Y(
        n368) );
  MX4X1 U1187 ( .A(n379), .B(n377), .C(n378), .D(n376), .S0(n3735), .S1(n3739), 
        .Y(n210) );
  MXI4X1 U1188 ( .A(\regfile[16][17] ), .B(\regfile[17][17] ), .C(
        \regfile[18][17] ), .D(\regfile[19][17] ), .S0(n3758), .S1(n3753), .Y(
        n379) );
  MXI4X1 U1189 ( .A(\regfile[24][17] ), .B(\regfile[25][17] ), .C(
        \regfile[26][17] ), .D(\regfile[27][17] ), .S0(n3758), .S1(n3751), .Y(
        n377) );
  MXI4X1 U1190 ( .A(\regfile[28][17] ), .B(\regfile[29][17] ), .C(
        \regfile[30][17] ), .D(\regfile[31][17] ), .S0(n3758), .S1(n3748), .Y(
        n376) );
  MX4X1 U1191 ( .A(n387), .B(n385), .C(n386), .D(n384), .S0(n3735), .S1(n3738), 
        .Y(n212) );
  MXI4X1 U1192 ( .A(\regfile[16][18] ), .B(\regfile[17][18] ), .C(
        \regfile[18][18] ), .D(\regfile[19][18] ), .S0(n3759), .S1(n3748), .Y(
        n387) );
  MXI4X1 U1193 ( .A(\regfile[24][18] ), .B(\regfile[25][18] ), .C(
        \regfile[26][18] ), .D(\regfile[27][18] ), .S0(n3759), .S1(n3754), .Y(
        n385) );
  MXI4X1 U1194 ( .A(\regfile[28][18] ), .B(\regfile[29][18] ), .C(
        \regfile[30][18] ), .D(\regfile[31][18] ), .S0(n3758), .S1(n3752), .Y(
        n384) );
  MX4X1 U1195 ( .A(n395), .B(n393), .C(n394), .D(n392), .S0(n3735), .S1(N19), 
        .Y(n214) );
  MXI4X1 U1196 ( .A(\regfile[16][19] ), .B(\regfile[17][19] ), .C(
        \regfile[18][19] ), .D(\regfile[19][19] ), .S0(n3759), .S1(n3754), .Y(
        n395) );
  MXI4X1 U1197 ( .A(\regfile[24][19] ), .B(\regfile[25][19] ), .C(
        \regfile[26][19] ), .D(\regfile[27][19] ), .S0(n3759), .S1(n3755), .Y(
        n393) );
  MXI4X1 U1198 ( .A(\regfile[28][19] ), .B(\regfile[29][19] ), .C(
        \regfile[30][19] ), .D(\regfile[31][19] ), .S0(n3759), .S1(n3743), .Y(
        n392) );
  MX4X1 U1199 ( .A(n403), .B(n401), .C(n402), .D(n400), .S0(n3736), .S1(n3740), 
        .Y(n216) );
  MXI4X1 U1200 ( .A(\regfile[16][20] ), .B(\regfile[17][20] ), .C(
        \regfile[18][20] ), .D(\regfile[19][20] ), .S0(n3760), .S1(n3753), .Y(
        n403) );
  MXI4X1 U1201 ( .A(\regfile[24][20] ), .B(\regfile[25][20] ), .C(
        \regfile[26][20] ), .D(\regfile[27][20] ), .S0(n3759), .S1(n3743), .Y(
        n401) );
  MXI4X1 U1202 ( .A(\regfile[28][20] ), .B(\regfile[29][20] ), .C(
        \regfile[30][20] ), .D(\regfile[31][20] ), .S0(n3759), .S1(n3742), .Y(
        n400) );
  MX4X1 U1203 ( .A(n411), .B(n409), .C(n410), .D(n408), .S0(n3736), .S1(n3740), 
        .Y(n218) );
  MXI4X1 U1204 ( .A(\regfile[16][21] ), .B(\regfile[17][21] ), .C(
        \regfile[18][21] ), .D(\regfile[19][21] ), .S0(n3760), .S1(n3746), .Y(
        n411) );
  MXI4X1 U1205 ( .A(\regfile[24][21] ), .B(\regfile[25][21] ), .C(
        \regfile[26][21] ), .D(\regfile[27][21] ), .S0(n3760), .S1(n3743), .Y(
        n409) );
  MXI4X1 U1206 ( .A(\regfile[28][21] ), .B(\regfile[29][21] ), .C(
        \regfile[30][21] ), .D(\regfile[31][21] ), .S0(n3760), .S1(n3748), .Y(
        n408) );
  MX4X1 U1207 ( .A(n419), .B(n417), .C(n418), .D(n416), .S0(n3736), .S1(N19), 
        .Y(n220) );
  MXI4X1 U1208 ( .A(\regfile[16][22] ), .B(\regfile[17][22] ), .C(
        \regfile[18][22] ), .D(\regfile[19][22] ), .S0(n3761), .S1(n3742), .Y(
        n419) );
  MXI4X1 U1209 ( .A(\regfile[24][22] ), .B(\regfile[25][22] ), .C(
        \regfile[26][22] ), .D(\regfile[27][22] ), .S0(n3760), .S1(n3751), .Y(
        n417) );
  MXI4X1 U1210 ( .A(\regfile[28][22] ), .B(\regfile[29][22] ), .C(
        \regfile[30][22] ), .D(\regfile[31][22] ), .S0(n3760), .S1(n3743), .Y(
        n416) );
  MX4X1 U1211 ( .A(n427), .B(n425), .C(n426), .D(n424), .S0(n3736), .S1(n3739), 
        .Y(n222) );
  MXI4X1 U1212 ( .A(\regfile[16][23] ), .B(\regfile[17][23] ), .C(
        \regfile[18][23] ), .D(\regfile[19][23] ), .S0(n3761), .S1(n3742), .Y(
        n427) );
  MXI4X1 U1213 ( .A(\regfile[24][23] ), .B(\regfile[25][23] ), .C(
        \regfile[26][23] ), .D(\regfile[27][23] ), .S0(n3761), .S1(n3743), .Y(
        n425) );
  MXI4X1 U1214 ( .A(\regfile[28][23] ), .B(\regfile[29][23] ), .C(
        \regfile[30][23] ), .D(\regfile[31][23] ), .S0(n3761), .S1(n3748), .Y(
        n424) );
  MX4X1 U1215 ( .A(n435), .B(n433), .C(n434), .D(n432), .S0(n3736), .S1(N19), 
        .Y(n225) );
  MXI4X1 U1216 ( .A(\regfile[16][24] ), .B(\regfile[17][24] ), .C(
        \regfile[18][24] ), .D(\regfile[19][24] ), .S0(n3762), .S1(n3751), .Y(
        n435) );
  MXI4X1 U1217 ( .A(\regfile[24][24] ), .B(\regfile[25][24] ), .C(
        \regfile[26][24] ), .D(\regfile[27][24] ), .S0(n3761), .S1(n3753), .Y(
        n433) );
  MXI4X1 U1218 ( .A(\regfile[28][24] ), .B(\regfile[29][24] ), .C(
        \regfile[30][24] ), .D(\regfile[31][24] ), .S0(n3761), .S1(n3742), .Y(
        n432) );
  MX4X1 U1219 ( .A(n443), .B(n441), .C(n442), .D(n440), .S0(n3736), .S1(N19), 
        .Y(n227) );
  MXI4X1 U1220 ( .A(\regfile[16][25] ), .B(\regfile[17][25] ), .C(
        \regfile[18][25] ), .D(\regfile[19][25] ), .S0(n3762), .S1(n3755), .Y(
        n443) );
  MXI4X1 U1221 ( .A(\regfile[24][25] ), .B(\regfile[25][25] ), .C(
        \regfile[26][25] ), .D(\regfile[27][25] ), .S0(n3762), .S1(n3747), .Y(
        n441) );
  MXI4X1 U1222 ( .A(\regfile[28][25] ), .B(\regfile[29][25] ), .C(
        \regfile[30][25] ), .D(\regfile[31][25] ), .S0(n3762), .S1(n3747), .Y(
        n440) );
  MX4X1 U1223 ( .A(n451), .B(n449), .C(n450), .D(n448), .S0(n3737), .S1(n3740), 
        .Y(n229) );
  MXI4X1 U1224 ( .A(\regfile[16][26] ), .B(\regfile[17][26] ), .C(
        \regfile[18][26] ), .D(\regfile[19][26] ), .S0(n3762), .S1(n3746), .Y(
        n451) );
  MXI4X1 U1225 ( .A(\regfile[24][26] ), .B(\regfile[25][26] ), .C(
        \regfile[26][26] ), .D(\regfile[27][26] ), .S0(n3762), .S1(n3742), .Y(
        n449) );
  MXI4X1 U1226 ( .A(\regfile[28][26] ), .B(\regfile[29][26] ), .C(
        \regfile[30][26] ), .D(\regfile[31][26] ), .S0(n3762), .S1(n3743), .Y(
        n448) );
  MX4X1 U1227 ( .A(n459), .B(n457), .C(n458), .D(n456), .S0(n3737), .S1(n3740), 
        .Y(n231) );
  MXI4X1 U1228 ( .A(\regfile[16][27] ), .B(\regfile[17][27] ), .C(
        \regfile[18][27] ), .D(\regfile[19][27] ), .S0(n3763), .S1(n3748), .Y(
        n459) );
  MXI4X1 U1229 ( .A(\regfile[24][27] ), .B(\regfile[25][27] ), .C(
        \regfile[26][27] ), .D(\regfile[27][27] ), .S0(n3763), .S1(n3755), .Y(
        n457) );
  MXI4X1 U1230 ( .A(\regfile[28][27] ), .B(\regfile[29][27] ), .C(
        \regfile[30][27] ), .D(\regfile[31][27] ), .S0(n3763), .S1(n3748), .Y(
        n456) );
  MX4X1 U1231 ( .A(n467), .B(n465), .C(n466), .D(n464), .S0(n3737), .S1(n3740), 
        .Y(n233) );
  MXI4X1 U1232 ( .A(\regfile[16][28] ), .B(\regfile[17][28] ), .C(
        \regfile[18][28] ), .D(\regfile[19][28] ), .S0(n3763), .S1(n3744), .Y(
        n467) );
  MXI4X1 U1233 ( .A(\regfile[24][28] ), .B(\regfile[25][28] ), .C(
        \regfile[26][28] ), .D(\regfile[27][28] ), .S0(n3763), .S1(n3742), .Y(
        n465) );
  MXI4X1 U1234 ( .A(\regfile[28][28] ), .B(\regfile[29][28] ), .C(
        \regfile[30][28] ), .D(\regfile[31][28] ), .S0(n3763), .S1(n3751), .Y(
        n464) );
  MX4X1 U1235 ( .A(n475), .B(n473), .C(n474), .D(n472), .S0(n3737), .S1(n3740), 
        .Y(n235) );
  MXI4X1 U1236 ( .A(\regfile[16][29] ), .B(\regfile[17][29] ), .C(
        \regfile[18][29] ), .D(\regfile[19][29] ), .S0(n3764), .S1(n3744), .Y(
        n475) );
  MXI4X1 U1237 ( .A(\regfile[24][29] ), .B(\regfile[25][29] ), .C(
        \regfile[26][29] ), .D(\regfile[27][29] ), .S0(n3764), .S1(n3744), .Y(
        n473) );
  MXI4X1 U1238 ( .A(\regfile[28][29] ), .B(\regfile[29][29] ), .C(
        \regfile[30][29] ), .D(\regfile[31][29] ), .S0(n3764), .S1(n3744), .Y(
        n472) );
  MX4X1 U1239 ( .A(n483), .B(n481), .C(n482), .D(n480), .S0(n3737), .S1(n3740), 
        .Y(n237) );
  MXI4X1 U1240 ( .A(\regfile[16][30] ), .B(\regfile[17][30] ), .C(
        \regfile[18][30] ), .D(\regfile[19][30] ), .S0(n3764), .S1(n3744), .Y(
        n483) );
  MXI4X1 U1241 ( .A(\regfile[24][30] ), .B(\regfile[25][30] ), .C(
        \regfile[26][30] ), .D(\regfile[27][30] ), .S0(n3764), .S1(n3744), .Y(
        n481) );
  MXI4X1 U1242 ( .A(\regfile[28][30] ), .B(\regfile[29][30] ), .C(
        \regfile[30][30] ), .D(\regfile[31][30] ), .S0(n3764), .S1(n3744), .Y(
        n480) );
  MX4X1 U1243 ( .A(n491), .B(n489), .C(n490), .D(n488), .S0(n3737), .S1(n3740), 
        .Y(n239) );
  MXI4X1 U1244 ( .A(\regfile[16][31] ), .B(\regfile[17][31] ), .C(
        \regfile[18][31] ), .D(\regfile[19][31] ), .S0(n3765), .S1(n3744), .Y(
        n491) );
  MXI4X1 U1245 ( .A(\regfile[24][31] ), .B(\regfile[25][31] ), .C(
        \regfile[26][31] ), .D(\regfile[27][31] ), .S0(n3765), .S1(n3744), .Y(
        n489) );
  MXI4X1 U1246 ( .A(\regfile[28][31] ), .B(\regfile[29][31] ), .C(
        \regfile[30][31] ), .D(\regfile[31][31] ), .S0(n3765), .S1(n3744), .Y(
        n488) );
  MX4X1 U1247 ( .A(n3844), .B(n3842), .C(n3843), .D(n3841), .S0(N25), .S1(
        n4265), .Y(n3778) );
  MXI4X1 U1248 ( .A(\regfile[16][0] ), .B(\regfile[17][0] ), .C(
        \regfile[18][0] ), .D(\regfile[19][0] ), .S0(n4290), .S1(n4277), .Y(
        n3844) );
  MXI4X1 U1249 ( .A(\regfile[24][0] ), .B(\regfile[25][0] ), .C(
        \regfile[26][0] ), .D(\regfile[27][0] ), .S0(n4290), .S1(n4270), .Y(
        n3842) );
  MXI4X1 U1250 ( .A(\regfile[28][0] ), .B(\regfile[29][0] ), .C(
        \regfile[30][0] ), .D(\regfile[31][0] ), .S0(n4290), .S1(n4277), .Y(
        n3841) );
  MX4X1 U1251 ( .A(n3852), .B(n3850), .C(n3851), .D(n3849), .S0(n4426), .S1(
        n4262), .Y(n3780) );
  MXI4X1 U1252 ( .A(\regfile[16][1] ), .B(\regfile[17][1] ), .C(
        \regfile[18][1] ), .D(\regfile[19][1] ), .S0(n4291), .S1(n4274), .Y(
        n3852) );
  MXI4X1 U1253 ( .A(\regfile[24][1] ), .B(\regfile[25][1] ), .C(
        \regfile[26][1] ), .D(\regfile[27][1] ), .S0(n4290), .S1(n4279), .Y(
        n3850) );
  MXI4X1 U1254 ( .A(\regfile[28][1] ), .B(\regfile[29][1] ), .C(
        \regfile[30][1] ), .D(\regfile[31][1] ), .S0(n4290), .S1(n4275), .Y(
        n3849) );
  MX4X1 U1255 ( .A(n243), .B(n241), .C(n242), .D(n240), .S0(n3733), .S1(n3739), 
        .Y(n157) );
  MXI4X1 U1256 ( .A(\regfile[16][0] ), .B(\regfile[17][0] ), .C(
        \regfile[18][0] ), .D(\regfile[19][0] ), .S0(n3765), .S1(n3745), .Y(
        n243) );
  MXI4X1 U1257 ( .A(\regfile[24][0] ), .B(\regfile[25][0] ), .C(
        \regfile[26][0] ), .D(\regfile[27][0] ), .S0(n3765), .S1(n3745), .Y(
        n241) );
  MXI4X1 U1258 ( .A(\regfile[28][0] ), .B(\regfile[29][0] ), .C(
        \regfile[30][0] ), .D(\regfile[31][0] ), .S0(n3765), .S1(n3745), .Y(
        n240) );
  MX4X1 U1259 ( .A(n251), .B(n249), .C(n250), .D(n248), .S0(n3734), .S1(n3740), 
        .Y(n159) );
  MXI4X1 U1260 ( .A(\regfile[16][1] ), .B(\regfile[17][1] ), .C(
        \regfile[18][1] ), .D(\regfile[19][1] ), .S0(n3766), .S1(n3745), .Y(
        n251) );
  MXI4X1 U1261 ( .A(\regfile[24][1] ), .B(\regfile[25][1] ), .C(
        \regfile[26][1] ), .D(\regfile[27][1] ), .S0(n3765), .S1(n3745), .Y(
        n249) );
  MXI4X1 U1262 ( .A(\regfile[28][1] ), .B(\regfile[29][1] ), .C(
        \regfile[30][1] ), .D(\regfile[31][1] ), .S0(n3765), .S1(n3745), .Y(
        n248) );
  MX4X1 U1264 ( .A(n3992), .B(n3990), .C(n3991), .D(n3989), .S0(N25), .S1(
        n4263), .Y(n3813) );
  MX4X1 U1265 ( .A(n4032), .B(n4030), .C(n4031), .D(n4029), .S0(n4261), .S1(
        n4264), .Y(n3823) );
  MX4X1 U1267 ( .A(n3856), .B(n3854), .C(n3855), .D(n3853), .S0(n4258), .S1(
        N24), .Y(n3779) );
  MX4X1 U1268 ( .A(n3864), .B(n3862), .C(n3863), .D(n3861), .S0(n4259), .S1(
        n4262), .Y(n3781) );
  MX4X1 U1269 ( .A(n3872), .B(n3870), .C(n3871), .D(n3869), .S0(n4259), .S1(
        n4262), .Y(n3783) );
  MX4X1 U1270 ( .A(n3888), .B(n3886), .C(n3887), .D(n3885), .S0(n4259), .S1(
        n4262), .Y(n3787) );
  MX4X1 U1271 ( .A(n3912), .B(n3910), .C(n3911), .D(n3909), .S0(N25), .S1(N24), 
        .Y(n3793) );
  MX4X1 U1272 ( .A(n3920), .B(n3918), .C(n3919), .D(n3917), .S0(N25), .S1(N24), 
        .Y(n3795) );
  MX4X1 U1275 ( .A(n3936), .B(n3934), .C(n3935), .D(n3933), .S0(n4258), .S1(
        N24), .Y(n3799) );
  MX4X1 U1278 ( .A(n3952), .B(n3950), .C(n3951), .D(n3949), .S0(n4258), .S1(
        N24), .Y(n3803) );
  MX4X1 U1280 ( .A(n3960), .B(n3958), .C(n3959), .D(n3957), .S0(N25), .S1(
        n4263), .Y(n3805) );
  MX4X1 U1282 ( .A(n3968), .B(n3966), .C(n3967), .D(n3965), .S0(N25), .S1(
        n4263), .Y(n3807) );
  MX4X1 U1288 ( .A(n4040), .B(n4038), .C(n4039), .D(n4037), .S0(n4261), .S1(
        n4264), .Y(n3825) );
  MX4X1 U1289 ( .A(n4048), .B(n4046), .C(n4047), .D(n4045), .S0(n4261), .S1(
        n4264), .Y(n3827) );
  MX4X1 U1291 ( .A(n4056), .B(n4054), .C(n4055), .D(n4053), .S0(N25), .S1(
        n4265), .Y(n3829) );
  MX4X1 U1293 ( .A(n4064), .B(n4062), .C(n4063), .D(n4061), .S0(N25), .S1(
        n4265), .Y(n3831) );
  MX4X1 U1295 ( .A(n4072), .B(n4070), .C(n4071), .D(n4069), .S0(N25), .S1(
        n4265), .Y(n3833) );
  MX4X1 U1296 ( .A(n4080), .B(n4078), .C(n4079), .D(n4077), .S0(N25), .S1(
        n4265), .Y(n3835) );
  MX4X1 U1298 ( .A(n4088), .B(n4086), .C(n4087), .D(n4085), .S0(N25), .S1(
        n4265), .Y(n3837) );
  NOR2BX1 U1301 ( .AN(n3750), .B(n92), .Y(n3727) );
  NOR2BX1 U1302 ( .AN(n3750), .B(\regfile[3][1] ), .Y(n3722) );
  NOR2BX1 U1303 ( .AN(n3750), .B(\regfile[3][2] ), .Y(n3717) );
  NOR2BX1 U1304 ( .AN(n3750), .B(\regfile[3][3] ), .Y(n3712) );
  NOR2BX1 U1305 ( .AN(n3750), .B(n90), .Y(n3707) );
  NOR2BX1 U1306 ( .AN(n3749), .B(\regfile[3][5] ), .Y(n3702) );
  NOR2BX1 U1307 ( .AN(n3750), .B(\regfile[3][6] ), .Y(n3697) );
  NOR2BX1 U1308 ( .AN(n3749), .B(n89), .Y(n3692) );
  NOR2BX1 U1309 ( .AN(n3749), .B(\regfile[3][8] ), .Y(n1777) );
  NOR2BX1 U1310 ( .AN(n3749), .B(\regfile[3][9] ), .Y(n1741) );
  NOR2BX1 U1311 ( .AN(n3749), .B(n88), .Y(n1731) );
  NOR2BX1 U1312 ( .AN(n3749), .B(\regfile[3][11] ), .Y(n1721) );
  NOR2BX1 U1313 ( .AN(n3750), .B(\regfile[3][12] ), .Y(n1711) );
  NOR2BX1 U1314 ( .AN(n3749), .B(\regfile[3][13] ), .Y(n1701) );
  NOR2BX1 U1315 ( .AN(n3749), .B(\regfile[3][14] ), .Y(n1691) );
  NOR2BX1 U1316 ( .AN(n3749), .B(\regfile[3][15] ), .Y(n1681) );
  NOR2BX1 U1317 ( .AN(n3749), .B(\regfile[3][16] ), .Y(n628) );
  NOR2BX1 U1318 ( .AN(n3749), .B(\regfile[3][17] ), .Y(n566) );
  NOR2BX1 U1319 ( .AN(n3749), .B(n91), .Y(n561) );
  NOR2BX1 U1320 ( .AN(n3749), .B(n94), .Y(n556) );
  NOR2BX1 U1321 ( .AN(n3749), .B(n85), .Y(n551) );
  NOR2BX1 U1322 ( .AN(n3749), .B(\regfile[3][21] ), .Y(n546) );
  NOR2BX1 U1323 ( .AN(n3749), .B(\regfile[3][22] ), .Y(n541) );
  NOR2BX1 U1324 ( .AN(n3749), .B(n87), .Y(n536) );
  NOR2BX1 U1325 ( .AN(n3749), .B(\regfile[3][24] ), .Y(n531) );
  NOR2BX1 U1326 ( .AN(n3750), .B(\regfile[3][25] ), .Y(n526) );
  NOR2BX1 U1327 ( .AN(n3750), .B(\regfile[3][26] ), .Y(n521) );
  NOR2BX1 U1328 ( .AN(n3750), .B(\regfile[3][27] ), .Y(n516) );
  NOR2BX1 U1329 ( .AN(n3750), .B(\regfile[3][28] ), .Y(n511) );
  NOR2BX1 U1330 ( .AN(n3750), .B(\regfile[3][29] ), .Y(n506) );
  NOR2BX1 U1331 ( .AN(n3750), .B(\regfile[3][30] ), .Y(n501) );
  NOR2BX1 U1332 ( .AN(n3750), .B(\regfile[3][31] ), .Y(n496) );
  NOR2X1 U1333 ( .A(n3750), .B(\regfile[1][4] ), .Y(n3709) );
  NOR2X1 U1334 ( .A(n3750), .B(\regfile[1][6] ), .Y(n3699) );
  NOR2X1 U1335 ( .A(\regfile[1][0] ), .B(n3743), .Y(n3729) );
  NOR2X1 U1336 ( .A(n3742), .B(\regfile[1][1] ), .Y(n3724) );
  NOR2X1 U1338 ( .A(n3748), .B(\regfile[1][3] ), .Y(n3714) );
  NOR2X1 U1339 ( .A(\regfile[1][5] ), .B(n3755), .Y(n3704) );
  NOR2X1 U1340 ( .A(n3746), .B(\regfile[1][7] ), .Y(n3694) );
  NOR2X1 U1342 ( .A(n3742), .B(\regfile[1][9] ), .Y(n1749) );
  NOR2X1 U1343 ( .A(n3751), .B(\regfile[1][10] ), .Y(n1735) );
  NOR2X1 U1344 ( .A(n3743), .B(\regfile[1][11] ), .Y(n1725) );
  NOR2X1 U1345 ( .A(n3748), .B(\regfile[1][12] ), .Y(n1715) );
  NOR2X1 U1346 ( .A(n3755), .B(\regfile[1][13] ), .Y(n1705) );
  NOR2X1 U1347 ( .A(n3751), .B(\regfile[1][14] ), .Y(n1695) );
  NOR2X1 U1348 ( .A(n3743), .B(\regfile[1][15] ), .Y(n1685) );
  NOR2X1 U1350 ( .A(n3748), .B(\regfile[1][17] ), .Y(n568) );
  NOR2X1 U1351 ( .A(n3742), .B(\regfile[1][18] ), .Y(n563) );
  NOR2X1 U1352 ( .A(n3746), .B(\regfile[1][19] ), .Y(n558) );
  NOR2X1 U1353 ( .A(n3748), .B(\regfile[1][20] ), .Y(n553) );
  NOR2X1 U1354 ( .A(n3754), .B(\regfile[1][21] ), .Y(n548) );
  NOR2X1 U1355 ( .A(n3751), .B(\regfile[1][22] ), .Y(n543) );
  NOR2X1 U1356 ( .A(n3755), .B(\regfile[1][23] ), .Y(n538) );
  NOR2X1 U1357 ( .A(\regfile[1][24] ), .B(n3742), .Y(n533) );
  NOR2X1 U1358 ( .A(n3743), .B(\regfile[1][25] ), .Y(n528) );
  NOR2X1 U1359 ( .A(\regfile[1][26] ), .B(n3746), .Y(n523) );
  NOR2X1 U1360 ( .A(n3743), .B(\regfile[1][27] ), .Y(n518) );
  NOR2X1 U1361 ( .A(n3742), .B(\regfile[1][28] ), .Y(n513) );
  NOR2X1 U1362 ( .A(n3752), .B(\regfile[1][29] ), .Y(n508) );
  NOR2X1 U1364 ( .A(n3754), .B(\regfile[1][31] ), .Y(n498) );
  NOR2X1 U1365 ( .A(n4249), .B(n4248), .Y(n4251) );
  NOR2X1 U1366 ( .A(n4276), .B(n4301), .Y(n4248) );
  NOR2X1 U1367 ( .A(n3724), .B(n3723), .Y(n3726) );
  NOR2X1 U1368 ( .A(n3754), .B(n3776), .Y(n3723) );
  NOR2X1 U1371 ( .A(n4270), .B(n4301), .Y(n4243) );
  NAND2X1 U1372 ( .A(n4241), .B(n4240), .Y(n3872) );
  NOR2X1 U1373 ( .A(n4239), .B(n4238), .Y(n4241) );
  MXI2X1 U1374 ( .A(n1577), .B(n4237), .S0(n4298), .Y(n4240) );
  NOR2X1 U1375 ( .A(n4278), .B(n4301), .Y(n4238) );
  NAND2X1 U1376 ( .A(n4236), .B(n4235), .Y(n3880) );
  NOR2X1 U1377 ( .A(n4234), .B(n4233), .Y(n4236) );
  NOR2X1 U1379 ( .A(n4277), .B(n4301), .Y(n4233) );
  NAND2X1 U1380 ( .A(n4231), .B(n4230), .Y(n3888) );
  NOR2X1 U1381 ( .A(n4229), .B(n4228), .Y(n4231) );
  NOR2X1 U1383 ( .A(n4280), .B(n4301), .Y(n4228) );
  NAND2X1 U1384 ( .A(n4225), .B(n4226), .Y(n3896) );
  NOR2X1 U1385 ( .A(n4224), .B(n4223), .Y(n4226) );
  NOR2X1 U1387 ( .A(n4268), .B(n4301), .Y(n4223) );
  NAND2X1 U1388 ( .A(n4221), .B(n4220), .Y(n3904) );
  NOR2X1 U1389 ( .A(n4219), .B(n4218), .Y(n4221) );
  NOR2X1 U1391 ( .A(n4277), .B(n4301), .Y(n4218) );
  NAND2X1 U1392 ( .A(n4216), .B(n4215), .Y(n3912) );
  NOR2X1 U1393 ( .A(n4214), .B(n4213), .Y(n4216) );
  NOR2X1 U1395 ( .A(n4276), .B(n4301), .Y(n4213) );
  NAND2X1 U1396 ( .A(n4211), .B(n4210), .Y(n3920) );
  NOR2X1 U1397 ( .A(n4209), .B(n4208), .Y(n4211) );
  NOR2X1 U1399 ( .A(n4274), .B(n4301), .Y(n4208) );
  NAND2X1 U1400 ( .A(n4206), .B(n4205), .Y(n3928) );
  MXI2X1 U1401 ( .A(n1570), .B(n4202), .S0(n4298), .Y(n4205) );
  NOR2X1 U1402 ( .A(n4270), .B(n4300), .Y(n4203) );
  NAND2X1 U1403 ( .A(n4201), .B(n4200), .Y(n3936) );
  NOR2X1 U1404 ( .A(n4199), .B(n4198), .Y(n4201) );
  NOR2X1 U1406 ( .A(n4276), .B(n4301), .Y(n4198) );
  NAND2X1 U1407 ( .A(n4196), .B(n4195), .Y(n3944) );
  NOR2X1 U1408 ( .A(n4194), .B(n4193), .Y(n4196) );
  MXI2X1 U1409 ( .A(n1568), .B(n4192), .S0(n4298), .Y(n4195) );
  NOR2X1 U1410 ( .A(n4277), .B(n4301), .Y(n4193) );
  NAND2X1 U1411 ( .A(n4191), .B(n4190), .Y(n3952) );
  NOR2X1 U1412 ( .A(n4189), .B(n4188), .Y(n4191) );
  NOR2X1 U1414 ( .A(n4279), .B(n4301), .Y(n4188) );
  NAND2X1 U1415 ( .A(n4186), .B(n4185), .Y(n3960) );
  NOR2X1 U1416 ( .A(n4184), .B(n4183), .Y(n4186) );
  MXI2X1 U1417 ( .A(n1566), .B(n4182), .S0(n4298), .Y(n4185) );
  NOR2X1 U1418 ( .A(n4268), .B(n4299), .Y(n4183) );
  NAND2X1 U1419 ( .A(n4181), .B(n4180), .Y(n3968) );
  NOR2X1 U1420 ( .A(n4179), .B(n4178), .Y(n4181) );
  MXI2X1 U1421 ( .A(n1565), .B(n4177), .S0(n4299), .Y(n4180) );
  NOR2X1 U1422 ( .A(n4268), .B(n4300), .Y(n4178) );
  NAND2X1 U1423 ( .A(n4176), .B(n4175), .Y(n3976) );
  NOR2X1 U1424 ( .A(n4174), .B(n4173), .Y(n4176) );
  NOR2X1 U1426 ( .A(n4275), .B(n4300), .Y(n4173) );
  NAND2X1 U1427 ( .A(n4171), .B(n4170), .Y(n3984) );
  NOR2X1 U1428 ( .A(n4169), .B(n4168), .Y(n4171) );
  MXI2X1 U1429 ( .A(n1563), .B(n4167), .S0(n4299), .Y(n4170) );
  NOR2X1 U1430 ( .A(n4277), .B(n4300), .Y(n4168) );
  NAND2X1 U1431 ( .A(n4166), .B(n4165), .Y(n3992) );
  NOR2X1 U1432 ( .A(n4164), .B(n4163), .Y(n4166) );
  NOR2X1 U1434 ( .A(n4276), .B(n4300), .Y(n4163) );
  NAND2X1 U1435 ( .A(n4161), .B(n4160), .Y(n4000) );
  NOR2X1 U1436 ( .A(n4159), .B(n4158), .Y(n4161) );
  NOR2X1 U1438 ( .A(n4279), .B(n4300), .Y(n4158) );
  NAND2X1 U1439 ( .A(n4156), .B(n4155), .Y(n4008) );
  NOR2X1 U1440 ( .A(n4154), .B(n4153), .Y(n4156) );
  MXI2X1 U1441 ( .A(n1560), .B(n4152), .S0(n4299), .Y(n4155) );
  NOR2X1 U1442 ( .A(n4278), .B(n4300), .Y(n4153) );
  NAND2X1 U1443 ( .A(n4151), .B(n4150), .Y(n4016) );
  NOR2X1 U1444 ( .A(n4149), .B(n4148), .Y(n4151) );
  MXI2X1 U1445 ( .A(n1559), .B(n4147), .S0(n4299), .Y(n4150) );
  NOR2X1 U1446 ( .A(n4274), .B(n4300), .Y(n4148) );
  NAND2X1 U1447 ( .A(n4146), .B(n4145), .Y(n4024) );
  NOR2X1 U1448 ( .A(n4144), .B(n4143), .Y(n4146) );
  MXI2X1 U1449 ( .A(n1558), .B(n4142), .S0(n4299), .Y(n4145) );
  NOR2X1 U1450 ( .A(n4274), .B(n4300), .Y(n4143) );
  NAND2X1 U1451 ( .A(n4141), .B(n4140), .Y(n4032) );
  NOR2X1 U1452 ( .A(n4139), .B(n4138), .Y(n4141) );
  MXI2X1 U1453 ( .A(n1557), .B(n4137), .S0(n4299), .Y(n4140) );
  NOR2X1 U1454 ( .A(n4279), .B(n4300), .Y(n4138) );
  NAND2X1 U1455 ( .A(n4136), .B(n4135), .Y(n4040) );
  NOR2X1 U1456 ( .A(n4134), .B(n4133), .Y(n4136) );
  NOR2X1 U1458 ( .A(n4278), .B(n4300), .Y(n4133) );
  NAND2X1 U1459 ( .A(n4126), .B(n4125), .Y(n4056) );
  NOR2X1 U1460 ( .A(n4124), .B(n4123), .Y(n4126) );
  MXI2X1 U1461 ( .A(n1554), .B(n4122), .S0(n4299), .Y(n4125) );
  NOR2X1 U1462 ( .A(n4278), .B(n4299), .Y(n4123) );
  NAND2X1 U1463 ( .A(n4110), .B(n4111), .Y(n4080) );
  NOR2X1 U1464 ( .A(n4109), .B(n4108), .Y(n4111) );
  NOR2X1 U1466 ( .A(n4278), .B(n4301), .Y(n4108) );
  NAND2X1 U1467 ( .A(n4101), .B(n4100), .Y(n4096) );
  NOR2X1 U1468 ( .A(n4099), .B(n4098), .Y(n4101) );
  MXI2X1 U1469 ( .A(n1549), .B(n4097), .S0(n4299), .Y(n4100) );
  NOR2X1 U1470 ( .A(n4270), .B(n4301), .Y(n4098) );
  NAND2X1 U1471 ( .A(n3721), .B(n3720), .Y(n263) );
  NOR2X1 U1472 ( .A(n3719), .B(n3718), .Y(n3721) );
  NOR2X1 U1474 ( .A(n3746), .B(n3776), .Y(n3718) );
  NAND2X1 U1475 ( .A(n3716), .B(n3715), .Y(n271) );
  NOR2X1 U1476 ( .A(n3714), .B(n3713), .Y(n3716) );
  MXI2X1 U1477 ( .A(n1577), .B(n3712), .S0(n3773), .Y(n3715) );
  NOR2X1 U1478 ( .A(n3746), .B(n3776), .Y(n3713) );
  NAND2X1 U1479 ( .A(n3711), .B(n3710), .Y(n279) );
  NOR2X1 U1480 ( .A(n3709), .B(n3708), .Y(n3711) );
  MXI2X1 U1481 ( .A(n1576), .B(n3707), .S0(n3773), .Y(n3710) );
  NOR2X1 U1482 ( .A(n3743), .B(n3776), .Y(n3708) );
  NAND2X1 U1483 ( .A(n3706), .B(n3705), .Y(n287) );
  NOR2X1 U1484 ( .A(n3704), .B(n3703), .Y(n3706) );
  NOR2X1 U1485 ( .A(n3750), .B(n3776), .Y(n3703) );
  NAND2X1 U1486 ( .A(n3701), .B(n3700), .Y(n295) );
  NOR2X1 U1487 ( .A(n3699), .B(n3698), .Y(n3701) );
  NOR2X1 U1489 ( .A(n3755), .B(n3776), .Y(n3698) );
  NAND2X1 U1490 ( .A(n3696), .B(n3695), .Y(n303) );
  NOR2X1 U1491 ( .A(n3694), .B(n3693), .Y(n3696) );
  MXI2X1 U1492 ( .A(n1573), .B(n3692), .S0(n3773), .Y(n3695) );
  NOR2X1 U1493 ( .A(n3748), .B(n3776), .Y(n3693) );
  NAND2X1 U1494 ( .A(n3691), .B(n1787), .Y(n311) );
  NOR2X1 U1495 ( .A(n1781), .B(n1779), .Y(n3691) );
  NOR2X1 U1497 ( .A(n3752), .B(n3775), .Y(n1779) );
  NAND2X1 U1498 ( .A(n1761), .B(n1755), .Y(n319) );
  NOR2X1 U1499 ( .A(n1749), .B(n1747), .Y(n1761) );
  NOR2X1 U1501 ( .A(n3754), .B(n3776), .Y(n1747) );
  NAND2X1 U1502 ( .A(n1739), .B(n1737), .Y(n327) );
  NOR2X1 U1503 ( .A(n1735), .B(n1733), .Y(n1739) );
  MXI2X1 U1504 ( .A(n1570), .B(n1731), .S0(n3773), .Y(n1737) );
  NOR2X1 U1505 ( .A(n3753), .B(n3775), .Y(n1733) );
  NAND2X1 U1506 ( .A(n1729), .B(n1727), .Y(n335) );
  NOR2X1 U1507 ( .A(n1725), .B(n1723), .Y(n1729) );
  MXI2X1 U1508 ( .A(n1569), .B(n1721), .S0(n3773), .Y(n1727) );
  NOR2X1 U1509 ( .A(n3753), .B(n3776), .Y(n1723) );
  NAND2X1 U1510 ( .A(n1719), .B(n1717), .Y(n343) );
  NOR2X1 U1511 ( .A(n1715), .B(n1713), .Y(n1719) );
  MXI2X1 U1512 ( .A(n1568), .B(n1711), .S0(n3773), .Y(n1717) );
  NOR2X1 U1513 ( .A(n3746), .B(n3775), .Y(n1713) );
  NAND2X1 U1514 ( .A(n1709), .B(n1707), .Y(n351) );
  NOR2X1 U1515 ( .A(n1705), .B(n1703), .Y(n1709) );
  NOR2X1 U1517 ( .A(n3748), .B(n3776), .Y(n1703) );
  NAND2X1 U1518 ( .A(n1699), .B(n1697), .Y(n359) );
  NOR2X1 U1519 ( .A(n1695), .B(n1693), .Y(n1699) );
  MXI2X1 U1520 ( .A(n1566), .B(n1691), .S0(n3773), .Y(n1697) );
  NOR2X1 U1521 ( .A(n3752), .B(n3773), .Y(n1693) );
  NAND2X1 U1522 ( .A(n1689), .B(n1687), .Y(n367) );
  NOR2X1 U1523 ( .A(n1685), .B(n1683), .Y(n1689) );
  MXI2X1 U1524 ( .A(n1565), .B(n1681), .S0(n3774), .Y(n1687) );
  NOR2X1 U1525 ( .A(n3748), .B(n3776), .Y(n1683) );
  NAND2X1 U1526 ( .A(n1679), .B(n1677), .Y(n375) );
  NOR2X1 U1527 ( .A(n630), .B(n629), .Y(n1679) );
  NOR2X1 U1529 ( .A(n3753), .B(n3775), .Y(n629) );
  NAND2X1 U1530 ( .A(n627), .B(n623), .Y(n383) );
  NOR2X1 U1531 ( .A(n568), .B(n567), .Y(n627) );
  MXI2X1 U1532 ( .A(n1563), .B(n566), .S0(n3774), .Y(n623) );
  NOR2X1 U1533 ( .A(n3743), .B(n3775), .Y(n567) );
  NAND2X1 U1534 ( .A(n565), .B(n564), .Y(n391) );
  NOR2X1 U1535 ( .A(n563), .B(n562), .Y(n565) );
  MXI2X1 U1536 ( .A(n1562), .B(n561), .S0(n3774), .Y(n564) );
  NOR2X1 U1537 ( .A(n3752), .B(n3776), .Y(n562) );
  NAND2X1 U1538 ( .A(n560), .B(n559), .Y(n399) );
  NOR2X1 U1539 ( .A(n558), .B(n557), .Y(n560) );
  MXI2X1 U1540 ( .A(n1561), .B(n556), .S0(n3774), .Y(n559) );
  NOR2X1 U1541 ( .A(n3748), .B(n3775), .Y(n557) );
  NAND2X1 U1542 ( .A(n555), .B(n554), .Y(n407) );
  NOR2X1 U1543 ( .A(n553), .B(n552), .Y(n555) );
  MXI2X1 U1544 ( .A(n1560), .B(n551), .S0(n3774), .Y(n554) );
  NOR2X1 U1545 ( .A(n3746), .B(n3775), .Y(n552) );
  NAND2X1 U1546 ( .A(n550), .B(n549), .Y(n415) );
  NOR2X1 U1547 ( .A(n548), .B(n547), .Y(n550) );
  MXI2X1 U1548 ( .A(n1559), .B(n546), .S0(n3774), .Y(n549) );
  NOR2X1 U1549 ( .A(n3742), .B(n3775), .Y(n547) );
  NAND2X1 U1550 ( .A(n545), .B(n544), .Y(n423) );
  NOR2X1 U1551 ( .A(n543), .B(n542), .Y(n545) );
  MXI2X1 U1552 ( .A(n1558), .B(n541), .S0(n3774), .Y(n544) );
  NOR2X1 U1553 ( .A(n3752), .B(n3775), .Y(n542) );
  NAND2X1 U1554 ( .A(n540), .B(n539), .Y(n431) );
  NOR2X1 U1555 ( .A(n538), .B(n537), .Y(n540) );
  MXI2X1 U1556 ( .A(n1557), .B(n536), .S0(n3774), .Y(n539) );
  NOR2X1 U1557 ( .A(n3753), .B(n3775), .Y(n537) );
  NAND2X1 U1558 ( .A(n535), .B(n534), .Y(n439) );
  NOR2X1 U1559 ( .A(n533), .B(n532), .Y(n535) );
  NOR2X1 U1561 ( .A(n3754), .B(n3775), .Y(n532) );
  NAND2X1 U1562 ( .A(n525), .B(n524), .Y(n455) );
  NOR2X1 U1563 ( .A(n522), .B(n523), .Y(n525) );
  NOR2X1 U1565 ( .A(n3748), .B(n3775), .Y(n522) );
  NAND2X1 U1566 ( .A(n510), .B(n509), .Y(n479) );
  NOR2X1 U1567 ( .A(n508), .B(n507), .Y(n510) );
  NOR2X1 U1569 ( .A(n3754), .B(n3776), .Y(n507) );
  NAND2X1 U1570 ( .A(n500), .B(n499), .Y(n495) );
  NOR2X1 U1571 ( .A(n498), .B(n497), .Y(n500) );
  MXI2X1 U1572 ( .A(n1549), .B(n496), .S0(n3774), .Y(n499) );
  NOR2X1 U1573 ( .A(n3746), .B(n3776), .Y(n497) );
  NAND2X1 U1574 ( .A(n4256), .B(n4255), .Y(n3848) );
  NOR2X1 U1575 ( .A(n4254), .B(n4253), .Y(n4256) );
  NOR2X1 U1577 ( .A(n4269), .B(n4301), .Y(n4253) );
  NAND2X1 U1578 ( .A(n4131), .B(n4130), .Y(n4048) );
  NOR2X1 U1579 ( .A(n4129), .B(n4128), .Y(n4131) );
  NOR2X1 U1581 ( .A(n4274), .B(n4284), .Y(n4128) );
  NAND2X1 U1582 ( .A(n4121), .B(n4120), .Y(n4064) );
  NOR2X1 U1583 ( .A(n4119), .B(n4118), .Y(n4121) );
  MXI2X1 U1584 ( .A(n1553), .B(n4117), .S0(n4300), .Y(n4120) );
  NOR2X1 U1585 ( .A(n4269), .B(n4301), .Y(n4118) );
  NAND2X1 U1586 ( .A(n4116), .B(n4115), .Y(n4072) );
  NOR2X1 U1587 ( .A(n4114), .B(n4113), .Y(n4116) );
  MXI2X1 U1588 ( .A(n1552), .B(n4112), .S0(n4300), .Y(n4115) );
  NOR2X1 U1589 ( .A(n4269), .B(n4301), .Y(n4113) );
  NAND2X1 U1590 ( .A(n4106), .B(n4105), .Y(n4088) );
  NOR2X1 U1591 ( .A(n4104), .B(n4103), .Y(n4106) );
  MXI2X1 U1592 ( .A(n1550), .B(n4102), .S0(n4300), .Y(n4105) );
  NOR2X1 U1593 ( .A(n4276), .B(n4301), .Y(n4103) );
  NAND2X1 U1594 ( .A(n3731), .B(n3730), .Y(n247) );
  NOR2X1 U1595 ( .A(n3729), .B(n3728), .Y(n3731) );
  NOR2X1 U1597 ( .A(n3750), .B(n3776), .Y(n3728) );
  NAND2X1 U1598 ( .A(n530), .B(n529), .Y(n447) );
  NOR2X1 U1599 ( .A(n528), .B(n527), .Y(n530) );
  MXI2X1 U1600 ( .A(n1555), .B(n526), .S0(n3775), .Y(n529) );
  NOR2X1 U1601 ( .A(n3755), .B(n3775), .Y(n527) );
  NAND2X1 U1602 ( .A(n520), .B(n519), .Y(n463) );
  NOR2X1 U1603 ( .A(n518), .B(n517), .Y(n520) );
  NOR2X1 U1605 ( .A(n3742), .B(n3774), .Y(n517) );
  NAND2X1 U1606 ( .A(n515), .B(n514), .Y(n471) );
  NOR2X1 U1607 ( .A(n513), .B(n512), .Y(n515) );
  MXI2X1 U1608 ( .A(n1552), .B(n511), .S0(n3775), .Y(n514) );
  NOR2X1 U1609 ( .A(n3743), .B(n3776), .Y(n512) );
  NAND2X1 U1610 ( .A(n505), .B(n504), .Y(n487) );
  NOR2X1 U1611 ( .A(n503), .B(n502), .Y(n505) );
  NOR2X1 U1613 ( .A(n3746), .B(n3776), .Y(n502) );
  MXI4X1 U1614 ( .A(\regfile[20][0] ), .B(\regfile[21][0] ), .C(
        \regfile[22][0] ), .D(\regfile[23][0] ), .S0(n4290), .S1(n4270), .Y(
        n3843) );
  MXI4X1 U1615 ( .A(\regfile[4][0] ), .B(\regfile[5][0] ), .C(\regfile[6][0] ), 
        .D(\regfile[7][0] ), .S0(n4290), .S1(n4269), .Y(n3847) );
  MXI4X1 U1616 ( .A(\regfile[20][1] ), .B(\regfile[21][1] ), .C(
        \regfile[22][1] ), .D(\regfile[23][1] ), .S0(n4291), .S1(n4280), .Y(
        n3851) );
  MXI4X1 U1617 ( .A(\regfile[4][1] ), .B(\regfile[5][1] ), .C(\regfile[6][1] ), 
        .D(\regfile[7][1] ), .S0(n4291), .S1(n4269), .Y(n3855) );
  MXI4X1 U1618 ( .A(\regfile[20][2] ), .B(\regfile[21][2] ), .C(
        \regfile[22][2] ), .D(\regfile[23][2] ), .S0(n4291), .S1(n4278), .Y(
        n3859) );
  MXI4X1 U1619 ( .A(\regfile[4][2] ), .B(\regfile[5][2] ), .C(\regfile[6][2] ), 
        .D(\regfile[7][2] ), .S0(n4291), .S1(n4269), .Y(n3863) );
  MXI4X1 U1620 ( .A(\regfile[20][3] ), .B(\regfile[21][3] ), .C(
        \regfile[22][3] ), .D(\regfile[23][3] ), .S0(n4291), .S1(n4271), .Y(
        n3867) );
  MXI4X1 U1621 ( .A(\regfile[4][3] ), .B(\regfile[5][3] ), .C(\regfile[6][3] ), 
        .D(\regfile[7][3] ), .S0(n4292), .S1(n4271), .Y(n3871) );
  MXI4X1 U1622 ( .A(\regfile[20][4] ), .B(\regfile[21][4] ), .C(
        \regfile[22][4] ), .D(\regfile[23][4] ), .S0(n4292), .S1(n4271), .Y(
        n3875) );
  MXI4X1 U1623 ( .A(\regfile[4][4] ), .B(\regfile[5][4] ), .C(\regfile[6][4] ), 
        .D(\regfile[7][4] ), .S0(n4292), .S1(n4271), .Y(n3879) );
  MXI4X1 U1624 ( .A(\regfile[20][5] ), .B(\regfile[21][5] ), .C(
        \regfile[22][5] ), .D(\regfile[23][5] ), .S0(n4292), .S1(n4271), .Y(
        n3883) );
  MXI4X1 U1625 ( .A(\regfile[4][5] ), .B(\regfile[5][5] ), .C(\regfile[6][5] ), 
        .D(\regfile[7][5] ), .S0(n4293), .S1(n4271), .Y(n3887) );
  MXI4X1 U1626 ( .A(\regfile[20][6] ), .B(\regfile[21][6] ), .C(
        \regfile[22][6] ), .D(\regfile[23][6] ), .S0(n4293), .S1(n4272), .Y(
        n3891) );
  MXI4X1 U1627 ( .A(\regfile[4][6] ), .B(\regfile[5][6] ), .C(\regfile[6][6] ), 
        .D(\regfile[7][6] ), .S0(n4293), .S1(n4272), .Y(n3895) );
  MXI4X1 U1628 ( .A(\regfile[20][7] ), .B(\regfile[21][7] ), .C(
        \regfile[22][7] ), .D(\regfile[23][7] ), .S0(n4293), .S1(n4272), .Y(
        n3899) );
  MXI4X1 U1629 ( .A(\regfile[4][7] ), .B(\regfile[5][7] ), .C(\regfile[6][7] ), 
        .D(\regfile[7][7] ), .S0(n4294), .S1(n4272), .Y(n3903) );
  MXI4X1 U1630 ( .A(\regfile[20][8] ), .B(\regfile[21][8] ), .C(
        \regfile[22][8] ), .D(\regfile[23][8] ), .S0(n4294), .S1(n4272), .Y(
        n3907) );
  MXI4X1 U1631 ( .A(\regfile[4][8] ), .B(\regfile[5][8] ), .C(\regfile[6][8] ), 
        .D(\regfile[7][8] ), .S0(n4294), .S1(n4272), .Y(n3911) );
  MXI4X1 U1632 ( .A(\regfile[20][9] ), .B(\regfile[21][9] ), .C(
        \regfile[22][9] ), .D(\regfile[23][9] ), .S0(n4294), .S1(n4273), .Y(
        n3915) );
  MXI4X1 U1633 ( .A(\regfile[4][9] ), .B(\regfile[5][9] ), .C(\regfile[6][9] ), 
        .D(\regfile[7][9] ), .S0(n4295), .S1(n4273), .Y(n3919) );
  MXI4X1 U1634 ( .A(\regfile[20][10] ), .B(\regfile[21][10] ), .C(
        \regfile[22][10] ), .D(\regfile[23][10] ), .S0(n4295), .S1(n4273), .Y(
        n3923) );
  MXI4X1 U1635 ( .A(\regfile[4][10] ), .B(\regfile[5][10] ), .C(
        \regfile[6][10] ), .D(\regfile[7][10] ), .S0(n4295), .S1(n4273), .Y(
        n3927) );
  MXI4X1 U1636 ( .A(\regfile[20][11] ), .B(\regfile[21][11] ), .C(
        \regfile[22][11] ), .D(\regfile[23][11] ), .S0(n4295), .S1(n4273), .Y(
        n3931) );
  MXI4X1 U1637 ( .A(\regfile[4][11] ), .B(\regfile[5][11] ), .C(
        \regfile[6][11] ), .D(\regfile[7][11] ), .S0(n4296), .S1(n4273), .Y(
        n3935) );
  MXI4X1 U1638 ( .A(\regfile[20][12] ), .B(\regfile[21][12] ), .C(
        \regfile[22][12] ), .D(\regfile[23][12] ), .S0(n4296), .S1(n4266), .Y(
        n3939) );
  MXI4X1 U1639 ( .A(\regfile[4][12] ), .B(\regfile[5][12] ), .C(
        \regfile[6][12] ), .D(\regfile[7][12] ), .S0(n4294), .S1(n4272), .Y(
        n3943) );
  MXI4X1 U1640 ( .A(\regfile[20][13] ), .B(\regfile[21][13] ), .C(
        \regfile[22][13] ), .D(\regfile[23][13] ), .S0(n4296), .S1(n4268), .Y(
        n3947) );
  MXI4X1 U1641 ( .A(\regfile[4][13] ), .B(\regfile[5][13] ), .C(
        \regfile[6][13] ), .D(\regfile[7][13] ), .S0(n4296), .S1(n4270), .Y(
        n3951) );
  MXI4X1 U1642 ( .A(\regfile[20][14] ), .B(\regfile[21][14] ), .C(
        \regfile[22][14] ), .D(\regfile[23][14] ), .S0(n4297), .S1(n4267), .Y(
        n3955) );
  MXI4X1 U1643 ( .A(\regfile[4][14] ), .B(\regfile[5][14] ), .C(
        \regfile[6][14] ), .D(\regfile[7][14] ), .S0(n4297), .S1(n4277), .Y(
        n3959) );
  MXI4X1 U1644 ( .A(\regfile[20][15] ), .B(\regfile[21][15] ), .C(
        \regfile[22][15] ), .D(\regfile[23][15] ), .S0(n4297), .S1(n4266), .Y(
        n3963) );
  MXI4X1 U1645 ( .A(\regfile[4][15] ), .B(\regfile[5][15] ), .C(
        \regfile[6][15] ), .D(\regfile[7][15] ), .S0(n4294), .S1(n4272), .Y(
        n3967) );
  MXI4X1 U1646 ( .A(\regfile[20][16] ), .B(\regfile[21][16] ), .C(
        \regfile[22][16] ), .D(\regfile[23][16] ), .S0(n4283), .S1(n4279), .Y(
        n3971) );
  MXI4X1 U1647 ( .A(\regfile[4][16] ), .B(\regfile[5][16] ), .C(
        \regfile[6][16] ), .D(\regfile[7][16] ), .S0(n4283), .S1(n4275), .Y(
        n3975) );
  MXI4X1 U1648 ( .A(\regfile[20][17] ), .B(\regfile[21][17] ), .C(
        \regfile[22][17] ), .D(\regfile[23][17] ), .S0(n4283), .S1(n4279), .Y(
        n3979) );
  MXI4X1 U1649 ( .A(\regfile[4][17] ), .B(\regfile[5][17] ), .C(
        \regfile[6][17] ), .D(\regfile[7][17] ), .S0(n4283), .S1(n4267), .Y(
        n3983) );
  MXI4X1 U1650 ( .A(\regfile[20][18] ), .B(\regfile[21][18] ), .C(
        \regfile[22][18] ), .D(\regfile[23][18] ), .S0(n4284), .S1(n4269), .Y(
        n3987) );
  MXI4X1 U1651 ( .A(\regfile[4][18] ), .B(\regfile[5][18] ), .C(
        \regfile[6][18] ), .D(\regfile[7][18] ), .S0(n4284), .S1(n4277), .Y(
        n3991) );
  MXI4X1 U1652 ( .A(\regfile[20][19] ), .B(\regfile[21][19] ), .C(
        \regfile[22][19] ), .D(\regfile[23][19] ), .S0(n4284), .S1(n4279), .Y(
        n3995) );
  MXI4X1 U1653 ( .A(\regfile[4][19] ), .B(\regfile[5][19] ), .C(
        \regfile[6][19] ), .D(\regfile[7][19] ), .S0(n4284), .S1(n4274), .Y(
        n3999) );
  MXI4X1 U1654 ( .A(\regfile[20][20] ), .B(\regfile[21][20] ), .C(
        \regfile[22][20] ), .D(\regfile[23][20] ), .S0(n4285), .S1(n4267), .Y(
        n4003) );
  MXI4X1 U1655 ( .A(\regfile[4][20] ), .B(\regfile[5][20] ), .C(
        \regfile[6][20] ), .D(\regfile[7][20] ), .S0(n4285), .S1(n4267), .Y(
        n4007) );
  MXI4X1 U1656 ( .A(\regfile[20][21] ), .B(\regfile[21][21] ), .C(
        \regfile[22][21] ), .D(\regfile[23][21] ), .S0(n4285), .S1(n4266), .Y(
        n4011) );
  MXI4X1 U1657 ( .A(\regfile[4][21] ), .B(\regfile[5][21] ), .C(
        \regfile[6][21] ), .D(\regfile[7][21] ), .S0(n4285), .S1(n4266), .Y(
        n4015) );
  MXI4X1 U1658 ( .A(\regfile[20][22] ), .B(\regfile[21][22] ), .C(
        \regfile[22][22] ), .D(\regfile[23][22] ), .S0(n4285), .S1(n4280), .Y(
        n4019) );
  MXI4X1 U1659 ( .A(\regfile[4][22] ), .B(\regfile[5][22] ), .C(
        \regfile[6][22] ), .D(\regfile[7][22] ), .S0(n4286), .S1(n4267), .Y(
        n4023) );
  MXI4X1 U1660 ( .A(\regfile[20][23] ), .B(\regfile[21][23] ), .C(
        \regfile[22][23] ), .D(\regfile[23][23] ), .S0(n4286), .S1(n4269), .Y(
        n4027) );
  MXI4X1 U1661 ( .A(\regfile[4][23] ), .B(\regfile[5][23] ), .C(
        \regfile[6][23] ), .D(\regfile[7][23] ), .S0(n4286), .S1(n4274), .Y(
        n4031) );
  MXI4X1 U1662 ( .A(\regfile[20][24] ), .B(\regfile[21][24] ), .C(
        \regfile[22][24] ), .D(\regfile[23][24] ), .S0(n4286), .S1(n4270), .Y(
        n4035) );
  MXI4X1 U1663 ( .A(\regfile[4][24] ), .B(\regfile[5][24] ), .C(
        \regfile[6][24] ), .D(\regfile[7][24] ), .S0(n4287), .S1(n4276), .Y(
        n4039) );
  MXI4X1 U1664 ( .A(\regfile[20][25] ), .B(\regfile[21][25] ), .C(
        \regfile[22][25] ), .D(\regfile[23][25] ), .S0(n4287), .S1(n4268), .Y(
        n4043) );
  MXI4X1 U1665 ( .A(\regfile[4][25] ), .B(\regfile[5][25] ), .C(
        \regfile[6][25] ), .D(\regfile[7][25] ), .S0(n4287), .S1(n4277), .Y(
        n4047) );
  MXI4X1 U1666 ( .A(\regfile[20][26] ), .B(\regfile[21][26] ), .C(
        \regfile[22][26] ), .D(\regfile[23][26] ), .S0(n4287), .S1(n4267), .Y(
        n4051) );
  MXI4X1 U1667 ( .A(\regfile[4][26] ), .B(\regfile[5][26] ), .C(
        \regfile[6][26] ), .D(\regfile[7][26] ), .S0(n4288), .S1(n4278), .Y(
        n4055) );
  MXI4X1 U1668 ( .A(\regfile[20][27] ), .B(\regfile[21][27] ), .C(
        \regfile[22][27] ), .D(\regfile[23][27] ), .S0(n4288), .S1(n4280), .Y(
        n4059) );
  MXI4X1 U1669 ( .A(\regfile[4][27] ), .B(\regfile[5][27] ), .C(
        \regfile[6][27] ), .D(\regfile[7][27] ), .S0(n4288), .S1(n4274), .Y(
        n4063) );
  MXI4X1 U1670 ( .A(\regfile[20][28] ), .B(\regfile[21][28] ), .C(
        \regfile[22][28] ), .D(\regfile[23][28] ), .S0(n4288), .S1(n4278), .Y(
        n4067) );
  MXI4X1 U1671 ( .A(\regfile[4][28] ), .B(\regfile[5][28] ), .C(
        \regfile[6][28] ), .D(\regfile[7][28] ), .S0(n4289), .S1(n4271), .Y(
        n4071) );
  MXI4X1 U1672 ( .A(\regfile[20][29] ), .B(\regfile[21][29] ), .C(
        \regfile[22][29] ), .D(\regfile[23][29] ), .S0(n4289), .S1(n4278), .Y(
        n4075) );
  MXI4X1 U1673 ( .A(\regfile[4][29] ), .B(\regfile[5][29] ), .C(
        \regfile[6][29] ), .D(\regfile[7][29] ), .S0(n4289), .S1(n4278), .Y(
        n4079) );
  MXI4X1 U1674 ( .A(\regfile[20][30] ), .B(\regfile[21][30] ), .C(
        \regfile[22][30] ), .D(\regfile[23][30] ), .S0(n4289), .S1(n4278), .Y(
        n4083) );
  MXI4X1 U1675 ( .A(\regfile[4][30] ), .B(\regfile[5][30] ), .C(
        \regfile[6][30] ), .D(\regfile[7][30] ), .S0(n4290), .S1(n4271), .Y(
        n4087) );
  MXI4X1 U1676 ( .A(\regfile[20][31] ), .B(\regfile[21][31] ), .C(
        \regfile[22][31] ), .D(\regfile[23][31] ), .S0(n4290), .S1(n4271), .Y(
        n4091) );
  MXI4X1 U1677 ( .A(\regfile[4][31] ), .B(\regfile[5][31] ), .C(
        \regfile[6][31] ), .D(\regfile[7][31] ), .S0(n4297), .S1(n4266), .Y(
        n4095) );
  MXI4X1 U1678 ( .A(\regfile[20][0] ), .B(\regfile[21][0] ), .C(
        \regfile[22][0] ), .D(\regfile[23][0] ), .S0(n3765), .S1(n3745), .Y(
        n242) );
  MXI4X1 U1679 ( .A(\regfile[4][0] ), .B(\regfile[5][0] ), .C(\regfile[6][0] ), 
        .D(\regfile[7][0] ), .S0(n3765), .S1(n3745), .Y(n246) );
  MXI4X1 U1680 ( .A(\regfile[20][1] ), .B(\regfile[21][1] ), .C(
        \regfile[22][1] ), .D(\regfile[23][1] ), .S0(n3766), .S1(n3745), .Y(
        n250) );
  MXI4X1 U1681 ( .A(\regfile[4][1] ), .B(\regfile[5][1] ), .C(\regfile[6][1] ), 
        .D(\regfile[7][1] ), .S0(n3766), .S1(n3745), .Y(n254) );
  MXI4X1 U1682 ( .A(\regfile[20][2] ), .B(\regfile[21][2] ), .C(
        \regfile[22][2] ), .D(\regfile[23][2] ), .S0(n3766), .S1(n3745), .Y(
        n258) );
  MXI4X1 U1683 ( .A(\regfile[4][2] ), .B(\regfile[5][2] ), .C(\regfile[6][2] ), 
        .D(\regfile[7][2] ), .S0(n3766), .S1(n3745), .Y(n262) );
  MXI4X1 U1684 ( .A(\regfile[20][3] ), .B(\regfile[21][3] ), .C(
        \regfile[22][3] ), .D(\regfile[23][3] ), .S0(n3766), .S1(n3742), .Y(
        n266) );
  MXI4X1 U1717 ( .A(\regfile[4][3] ), .B(\regfile[5][3] ), .C(\regfile[6][3] ), 
        .D(\regfile[7][3] ), .S0(n3767), .S1(n3743), .Y(n270) );
  MXI4X1 U1718 ( .A(\regfile[20][4] ), .B(\regfile[21][4] ), .C(
        \regfile[22][4] ), .D(\regfile[23][4] ), .S0(n3767), .S1(n3746), .Y(
        n274) );
  MXI4X1 U1719 ( .A(\regfile[4][4] ), .B(\regfile[5][4] ), .C(\regfile[6][4] ), 
        .D(\regfile[7][4] ), .S0(n3767), .S1(n3755), .Y(n278) );
  MXI4X1 U1720 ( .A(\regfile[20][5] ), .B(\regfile[21][5] ), .C(
        \regfile[22][5] ), .D(\regfile[23][5] ), .S0(n3767), .S1(n3754), .Y(
        n282) );
  MXI4X1 U1721 ( .A(\regfile[4][5] ), .B(\regfile[5][5] ), .C(\regfile[6][5] ), 
        .D(\regfile[7][5] ), .S0(n3768), .S1(n3753), .Y(n286) );
  MXI4X1 U1722 ( .A(\regfile[20][6] ), .B(\regfile[21][6] ), .C(
        \regfile[22][6] ), .D(\regfile[23][6] ), .S0(n3768), .S1(n3745), .Y(
        n290) );
  MXI4X1 U1723 ( .A(\regfile[20][7] ), .B(\regfile[21][7] ), .C(
        \regfile[22][7] ), .D(\regfile[23][7] ), .S0(n3768), .S1(n3742), .Y(
        n298) );
  MXI4X1 U1724 ( .A(\regfile[20][8] ), .B(\regfile[21][8] ), .C(
        \regfile[22][8] ), .D(\regfile[23][8] ), .S0(n3769), .S1(n3751), .Y(
        n306) );
  MXI4X1 U1725 ( .A(\regfile[4][8] ), .B(\regfile[5][8] ), .C(\regfile[6][8] ), 
        .D(\regfile[7][8] ), .S0(n3769), .S1(n3745), .Y(n310) );
  MXI4X1 U1726 ( .A(\regfile[20][9] ), .B(\regfile[21][9] ), .C(
        \regfile[22][9] ), .D(\regfile[23][9] ), .S0(n3769), .S1(n3747), .Y(
        n314) );
  MXI4X1 U1727 ( .A(\regfile[4][9] ), .B(\regfile[5][9] ), .C(\regfile[6][9] ), 
        .D(\regfile[7][9] ), .S0(n3770), .S1(n3747), .Y(n318) );
  MXI4X1 U1728 ( .A(\regfile[20][10] ), .B(\regfile[21][10] ), .C(
        \regfile[22][10] ), .D(\regfile[23][10] ), .S0(n3770), .S1(n3747), .Y(
        n322) );
  MXI4X1 U1729 ( .A(\regfile[4][10] ), .B(\regfile[5][10] ), .C(
        \regfile[6][10] ), .D(\regfile[7][10] ), .S0(n3770), .S1(n3747), .Y(
        n326) );
  MXI4X1 U1730 ( .A(\regfile[20][11] ), .B(\regfile[21][11] ), .C(
        \regfile[22][11] ), .D(\regfile[23][11] ), .S0(n3770), .S1(n3747), .Y(
        n330) );
  MXI4X1 U1731 ( .A(\regfile[4][11] ), .B(\regfile[5][11] ), .C(
        \regfile[6][11] ), .D(\regfile[7][11] ), .S0(n3771), .S1(n3747), .Y(
        n334) );
  MXI4X1 U1732 ( .A(\regfile[20][12] ), .B(\regfile[21][12] ), .C(
        \regfile[22][12] ), .D(\regfile[23][12] ), .S0(n3771), .S1(n3746), .Y(
        n338) );
  MXI4X1 U1733 ( .A(\regfile[4][12] ), .B(\regfile[5][12] ), .C(
        \regfile[6][12] ), .D(\regfile[7][12] ), .S0(n3769), .S1(n3741), .Y(
        n342) );
  MXI4X1 U1734 ( .A(\regfile[20][13] ), .B(\regfile[21][13] ), .C(
        \regfile[22][13] ), .D(\regfile[23][13] ), .S0(n3771), .S1(n3742), .Y(
        n346) );
  MXI4X1 U1735 ( .A(\regfile[4][13] ), .B(\regfile[5][13] ), .C(
        \regfile[6][13] ), .D(\regfile[7][13] ), .S0(n3771), .S1(n3753), .Y(
        n350) );
  MXI4X1 U1736 ( .A(\regfile[20][14] ), .B(\regfile[21][14] ), .C(
        \regfile[22][14] ), .D(\regfile[23][14] ), .S0(n3772), .S1(n3754), .Y(
        n354) );
  MXI4X1 U1737 ( .A(\regfile[4][14] ), .B(\regfile[5][14] ), .C(
        \regfile[6][14] ), .D(\regfile[7][14] ), .S0(n3772), .S1(n3755), .Y(
        n358) );
  MXI4X1 U1738 ( .A(\regfile[20][15] ), .B(\regfile[21][15] ), .C(
        \regfile[22][15] ), .D(\regfile[23][15] ), .S0(n3772), .S1(n3752), .Y(
        n362) );
  MXI4X1 U1739 ( .A(\regfile[4][15] ), .B(\regfile[5][15] ), .C(
        \regfile[6][15] ), .D(\regfile[7][15] ), .S0(n3769), .S1(n3753), .Y(
        n366) );
  MXI4X1 U1740 ( .A(\regfile[20][16] ), .B(\regfile[21][16] ), .C(
        \regfile[22][16] ), .D(\regfile[23][16] ), .S0(n3758), .S1(n3743), .Y(
        n370) );
  MXI4X1 U1741 ( .A(\regfile[4][16] ), .B(\regfile[5][16] ), .C(
        \regfile[6][16] ), .D(\regfile[7][16] ), .S0(n3758), .S1(n3754), .Y(
        n374) );
  MXI4X1 U1742 ( .A(\regfile[20][17] ), .B(\regfile[21][17] ), .C(
        \regfile[22][17] ), .D(\regfile[23][17] ), .S0(n3758), .S1(n3742), .Y(
        n378) );
  MXI4X1 U1743 ( .A(\regfile[4][17] ), .B(\regfile[5][17] ), .C(
        \regfile[6][17] ), .D(\regfile[7][17] ), .S0(n3758), .S1(n3751), .Y(
        n382) );
  MXI4X1 U1744 ( .A(\regfile[20][18] ), .B(\regfile[21][18] ), .C(
        \regfile[22][18] ), .D(\regfile[23][18] ), .S0(n3759), .S1(n3753), .Y(
        n386) );
  MXI4X1 U1745 ( .A(\regfile[4][18] ), .B(\regfile[5][18] ), .C(
        \regfile[6][18] ), .D(\regfile[7][18] ), .S0(n3759), .S1(n3754), .Y(
        n390) );
  MXI4X1 U1746 ( .A(\regfile[20][19] ), .B(\regfile[21][19] ), .C(
        \regfile[22][19] ), .D(\regfile[23][19] ), .S0(n3759), .S1(n3748), .Y(
        n394) );
  MXI4X1 U1747 ( .A(\regfile[4][19] ), .B(\regfile[5][19] ), .C(
        \regfile[6][19] ), .D(\regfile[7][19] ), .S0(n3759), .S1(n3746), .Y(
        n398) );
  MXI4X1 U1748 ( .A(\regfile[20][20] ), .B(\regfile[21][20] ), .C(
        \regfile[22][20] ), .D(\regfile[23][20] ), .S0(n3760), .S1(n3755), .Y(
        n402) );
  MXI4X1 U1749 ( .A(\regfile[4][20] ), .B(\regfile[5][20] ), .C(
        \regfile[6][20] ), .D(\regfile[7][20] ), .S0(n3760), .S1(n3743), .Y(
        n406) );
  MXI4X1 U1752 ( .A(\regfile[20][21] ), .B(\regfile[21][21] ), .C(
        \regfile[22][21] ), .D(\regfile[23][21] ), .S0(n3760), .S1(n3742), .Y(
        n410) );
  MXI4X1 U1753 ( .A(\regfile[4][21] ), .B(\regfile[5][21] ), .C(
        \regfile[6][21] ), .D(\regfile[7][21] ), .S0(n3760), .S1(n3754), .Y(
        n414) );
  MXI4X1 U1756 ( .A(\regfile[20][22] ), .B(\regfile[21][22] ), .C(
        \regfile[22][22] ), .D(\regfile[23][22] ), .S0(n3760), .S1(n3744), .Y(
        n418) );
  MXI4X1 U1759 ( .A(\regfile[4][22] ), .B(\regfile[5][22] ), .C(
        \regfile[6][22] ), .D(\regfile[7][22] ), .S0(n3761), .S1(n3752), .Y(
        n422) );
  MXI4X1 U1767 ( .A(\regfile[20][23] ), .B(\regfile[21][23] ), .C(
        \regfile[22][23] ), .D(\regfile[23][23] ), .S0(n3761), .S1(n3748), .Y(
        n426) );
  MXI4X1 U1768 ( .A(\regfile[4][23] ), .B(\regfile[5][23] ), .C(
        \regfile[6][23] ), .D(\regfile[7][23] ), .S0(n3761), .S1(n3752), .Y(
        n430) );
  MXI4X1 U1769 ( .A(\regfile[20][24] ), .B(\regfile[21][24] ), .C(
        \regfile[22][24] ), .D(\regfile[23][24] ), .S0(n3761), .S1(n3742), .Y(
        n434) );
  MXI4X1 U1772 ( .A(\regfile[4][24] ), .B(\regfile[5][24] ), .C(
        \regfile[6][24] ), .D(\regfile[7][24] ), .S0(n3762), .S1(n3747), .Y(
        n438) );
  MXI4X1 U2678 ( .A(\regfile[20][25] ), .B(\regfile[21][25] ), .C(
        \regfile[22][25] ), .D(\regfile[23][25] ), .S0(n3762), .S1(n3751), .Y(
        n442) );
  MXI4X1 U2679 ( .A(\regfile[4][25] ), .B(\regfile[5][25] ), .C(
        \regfile[6][25] ), .D(\regfile[7][25] ), .S0(n3762), .S1(n3752), .Y(
        n446) );
  MXI4X1 U2680 ( .A(\regfile[20][26] ), .B(\regfile[21][26] ), .C(
        \regfile[22][26] ), .D(\regfile[23][26] ), .S0(n3762), .S1(n3751), .Y(
        n450) );
  MXI4X1 U2681 ( .A(\regfile[4][26] ), .B(\regfile[5][26] ), .C(
        \regfile[6][26] ), .D(\regfile[7][26] ), .S0(n3763), .S1(n3752), .Y(
        n454) );
  MXI4X1 U2682 ( .A(\regfile[20][27] ), .B(\regfile[21][27] ), .C(
        \regfile[22][27] ), .D(\regfile[23][27] ), .S0(n3763), .S1(n3748), .Y(
        n458) );
  MXI4X1 U2683 ( .A(\regfile[4][27] ), .B(\regfile[5][27] ), .C(
        \regfile[6][27] ), .D(\regfile[7][27] ), .S0(n3763), .S1(n3745), .Y(
        n462) );
  MXI4X1 U2684 ( .A(\regfile[20][28] ), .B(\regfile[21][28] ), .C(
        \regfile[22][28] ), .D(\regfile[23][28] ), .S0(n3763), .S1(n3746), .Y(
        n466) );
  MXI4X1 U2685 ( .A(\regfile[4][28] ), .B(\regfile[5][28] ), .C(
        \regfile[6][28] ), .D(\regfile[7][28] ), .S0(n3764), .S1(n3744), .Y(
        n470) );
  MXI4X1 U2686 ( .A(\regfile[20][29] ), .B(\regfile[21][29] ), .C(
        \regfile[22][29] ), .D(\regfile[23][29] ), .S0(n3764), .S1(n3744), .Y(
        n474) );
  MXI4X1 U2687 ( .A(\regfile[4][29] ), .B(\regfile[5][29] ), .C(
        \regfile[6][29] ), .D(\regfile[7][29] ), .S0(n3764), .S1(n3744), .Y(
        n478) );
  MXI4X1 U2688 ( .A(\regfile[20][30] ), .B(\regfile[21][30] ), .C(
        \regfile[22][30] ), .D(\regfile[23][30] ), .S0(n3764), .S1(n3744), .Y(
        n482) );
  MXI4X1 U2689 ( .A(\regfile[4][30] ), .B(\regfile[5][30] ), .C(
        \regfile[6][30] ), .D(\regfile[7][30] ), .S0(n3765), .S1(n3744), .Y(
        n486) );
  MXI4X1 U2690 ( .A(\regfile[20][31] ), .B(\regfile[21][31] ), .C(
        \regfile[22][31] ), .D(\regfile[23][31] ), .S0(n3765), .S1(n3744), .Y(
        n490) );
  MXI4X1 U2691 ( .A(\regfile[4][31] ), .B(\regfile[5][31] ), .C(
        \regfile[6][31] ), .D(\regfile[7][31] ), .S0(n3772), .S1(n3749), .Y(
        n494) );
  MXI4X1 U2692 ( .A(\regfile[12][0] ), .B(\regfile[13][0] ), .C(
        \regfile[14][0] ), .D(\regfile[15][0] ), .S0(n4290), .S1(n4275), .Y(
        n3845) );
  MXI4X1 U2693 ( .A(\regfile[12][1] ), .B(\regfile[13][1] ), .C(
        \regfile[14][1] ), .D(\regfile[15][1] ), .S0(n4291), .S1(n4276), .Y(
        n3853) );
  MXI4X1 U2694 ( .A(\regfile[12][2] ), .B(\regfile[13][2] ), .C(
        \regfile[14][2] ), .D(\regfile[15][2] ), .S0(n4291), .S1(n4268), .Y(
        n3861) );
  MXI4X1 U2695 ( .A(\regfile[12][3] ), .B(\regfile[13][3] ), .C(
        \regfile[14][3] ), .D(\regfile[15][3] ), .S0(n4292), .S1(n4271), .Y(
        n3869) );
  MXI4X1 U2696 ( .A(\regfile[12][4] ), .B(\regfile[13][4] ), .C(
        \regfile[14][4] ), .D(\regfile[15][4] ), .S0(n4292), .S1(n4271), .Y(
        n3877) );
  MXI4X1 U2697 ( .A(\regfile[12][5] ), .B(\regfile[13][5] ), .C(
        \regfile[14][5] ), .D(\regfile[15][5] ), .S0(n4293), .S1(n4271), .Y(
        n3885) );
  MXI4X1 U2698 ( .A(\regfile[12][6] ), .B(\regfile[13][6] ), .C(
        \regfile[14][6] ), .D(\regfile[15][6] ), .S0(n4293), .S1(n4272), .Y(
        n3893) );
  MXI4X1 U2699 ( .A(\regfile[12][7] ), .B(\regfile[13][7] ), .C(
        \regfile[14][7] ), .D(\regfile[15][7] ), .S0(n4293), .S1(n4272), .Y(
        n3901) );
  MXI4X1 U2700 ( .A(\regfile[12][8] ), .B(\regfile[13][8] ), .C(
        \regfile[14][8] ), .D(\regfile[15][8] ), .S0(n4294), .S1(n4272), .Y(
        n3909) );
  MXI4X1 U2701 ( .A(\regfile[12][9] ), .B(\regfile[13][9] ), .C(
        \regfile[14][9] ), .D(\regfile[15][9] ), .S0(n4294), .S1(n4273), .Y(
        n3917) );
  MXI4X1 U2702 ( .A(\regfile[12][10] ), .B(\regfile[13][10] ), .C(
        \regfile[14][10] ), .D(\regfile[15][10] ), .S0(n4295), .S1(n4273), .Y(
        n3925) );
  MXI4X1 U2703 ( .A(\regfile[12][11] ), .B(\regfile[13][11] ), .C(
        \regfile[14][11] ), .D(\regfile[15][11] ), .S0(n4295), .S1(n4273), .Y(
        n3933) );
  MXI4X1 U2704 ( .A(\regfile[12][12] ), .B(\regfile[13][12] ), .C(
        \regfile[14][12] ), .D(\regfile[15][12] ), .S0(n4296), .S1(n4266), .Y(
        n3941) );
  MXI4X1 U2705 ( .A(\regfile[12][13] ), .B(\regfile[13][13] ), .C(
        \regfile[14][13] ), .D(\regfile[15][13] ), .S0(n4296), .S1(n4272), .Y(
        n3949) );
  MXI4X1 U2706 ( .A(\regfile[12][14] ), .B(\regfile[13][14] ), .C(
        \regfile[14][14] ), .D(\regfile[15][14] ), .S0(n4297), .S1(n4273), .Y(
        n3957) );
  MXI4X1 U2707 ( .A(\regfile[12][15] ), .B(\regfile[13][15] ), .C(
        \regfile[14][15] ), .D(\regfile[15][15] ), .S0(n4297), .S1(n4279), .Y(
        n3965) );
  MXI4X1 U2708 ( .A(\regfile[12][16] ), .B(\regfile[13][16] ), .C(
        \regfile[14][16] ), .D(\regfile[15][16] ), .S0(n4283), .S1(n4270), .Y(
        n3973) );
  MXI4X1 U2709 ( .A(\regfile[12][17] ), .B(\regfile[13][17] ), .C(
        \regfile[14][17] ), .D(\regfile[15][17] ), .S0(n4283), .S1(n4267), .Y(
        n3981) );
  MXI4X1 U2710 ( .A(\regfile[12][18] ), .B(\regfile[13][18] ), .C(
        \regfile[14][18] ), .D(\regfile[15][18] ), .S0(n4284), .S1(n4268), .Y(
        n3989) );
  MXI4X1 U2711 ( .A(\regfile[12][19] ), .B(\regfile[13][19] ), .C(
        \regfile[14][19] ), .D(\regfile[15][19] ), .S0(n4284), .S1(n4277), .Y(
        n3997) );
  MXI4X1 U2712 ( .A(\regfile[12][20] ), .B(\regfile[13][20] ), .C(
        \regfile[14][20] ), .D(\regfile[15][20] ), .S0(n4285), .S1(n4267), .Y(
        n4005) );
  MXI4X1 U2713 ( .A(\regfile[12][21] ), .B(\regfile[13][21] ), .C(
        \regfile[14][21] ), .D(\regfile[15][21] ), .S0(n4285), .S1(n4266), .Y(
        n4013) );
  MXI4X1 U2714 ( .A(\regfile[12][22] ), .B(\regfile[13][22] ), .C(
        \regfile[14][22] ), .D(\regfile[15][22] ), .S0(n4286), .S1(n4267), .Y(
        n4021) );
  MXI4X1 U2715 ( .A(\regfile[12][23] ), .B(\regfile[13][23] ), .C(
        \regfile[14][23] ), .D(\regfile[15][23] ), .S0(n4286), .S1(n4278), .Y(
        n4029) );
  MXI4X1 U2716 ( .A(\regfile[12][24] ), .B(\regfile[13][24] ), .C(
        \regfile[14][24] ), .D(\regfile[15][24] ), .S0(n4287), .S1(n4274), .Y(
        n4037) );
  MXI4X1 U2717 ( .A(\regfile[12][25] ), .B(\regfile[13][25] ), .C(
        \regfile[14][25] ), .D(\regfile[15][25] ), .S0(n4287), .S1(n4270), .Y(
        n4045) );
  MXI4X1 U2718 ( .A(\regfile[12][26] ), .B(\regfile[13][26] ), .C(
        \regfile[14][26] ), .D(\regfile[15][26] ), .S0(n4288), .S1(n4275), .Y(
        n4053) );
  MXI4X1 U2719 ( .A(\regfile[12][27] ), .B(\regfile[13][27] ), .C(
        \regfile[14][27] ), .D(\regfile[15][27] ), .S0(n4288), .S1(n4278), .Y(
        n4061) );
  MXI4X1 U2720 ( .A(\regfile[12][28] ), .B(\regfile[13][28] ), .C(
        \regfile[14][28] ), .D(\regfile[15][28] ), .S0(n4288), .S1(n4279), .Y(
        n4069) );
  MXI4X1 U2721 ( .A(\regfile[12][29] ), .B(\regfile[13][29] ), .C(
        \regfile[14][29] ), .D(\regfile[15][29] ), .S0(n4289), .S1(n4279), .Y(
        n4077) );
  MXI4X1 U2722 ( .A(\regfile[12][30] ), .B(\regfile[13][30] ), .C(
        \regfile[14][30] ), .D(\regfile[15][30] ), .S0(n4289), .S1(n4274), .Y(
        n4085) );
  MXI4X1 U2723 ( .A(\regfile[12][31] ), .B(\regfile[13][31] ), .C(
        \regfile[14][31] ), .D(\regfile[15][31] ), .S0(n4290), .S1(n4266), .Y(
        n4093) );
  MXI4X1 U2724 ( .A(\regfile[12][0] ), .B(\regfile[13][0] ), .C(
        \regfile[14][0] ), .D(\regfile[15][0] ), .S0(n3765), .S1(n3745), .Y(
        n244) );
  MXI4X1 U2725 ( .A(\regfile[12][1] ), .B(\regfile[13][1] ), .C(
        \regfile[14][1] ), .D(\regfile[15][1] ), .S0(n3766), .S1(n3745), .Y(
        n252) );
  MXI4X1 U2726 ( .A(\regfile[12][2] ), .B(\regfile[13][2] ), .C(
        \regfile[14][2] ), .D(\regfile[15][2] ), .S0(n3766), .S1(n3745), .Y(
        n260) );
  MXI4X1 U2727 ( .A(\regfile[12][3] ), .B(\regfile[13][3] ), .C(
        \regfile[14][3] ), .D(\regfile[15][3] ), .S0(n3767), .S1(n3754), .Y(
        n268) );
  MXI4X1 U2728 ( .A(\regfile[12][4] ), .B(\regfile[13][4] ), .C(
        \regfile[14][4] ), .D(\regfile[15][4] ), .S0(n3767), .S1(n3743), .Y(
        n276) );
  MXI4X1 U2729 ( .A(\regfile[12][5] ), .B(\regfile[13][5] ), .C(
        \regfile[14][5] ), .D(\regfile[15][5] ), .S0(n3768), .S1(n3751), .Y(
        n284) );
  MXI4X1 U2730 ( .A(\regfile[12][8] ), .B(\regfile[13][8] ), .C(
        \regfile[14][8] ), .D(\regfile[15][8] ), .S0(n3769), .S1(n3751), .Y(
        n308) );
  MXI4X1 U2731 ( .A(\regfile[12][9] ), .B(\regfile[13][9] ), .C(
        \regfile[14][9] ), .D(\regfile[15][9] ), .S0(n3769), .S1(n3747), .Y(
        n316) );
  MXI4X1 U2732 ( .A(\regfile[12][10] ), .B(\regfile[13][10] ), .C(
        \regfile[14][10] ), .D(\regfile[15][10] ), .S0(n3770), .S1(n3747), .Y(
        n324) );
  MXI4X1 U2733 ( .A(\regfile[12][11] ), .B(\regfile[13][11] ), .C(
        \regfile[14][11] ), .D(\regfile[15][11] ), .S0(n3770), .S1(n3747), .Y(
        n332) );
  MXI4X1 U2734 ( .A(\regfile[12][12] ), .B(\regfile[13][12] ), .C(
        \regfile[14][12] ), .D(\regfile[15][12] ), .S0(n3771), .S1(n3743), .Y(
        n340) );
  MXI4X1 U2735 ( .A(\regfile[12][13] ), .B(\regfile[13][13] ), .C(
        \regfile[14][13] ), .D(\regfile[15][13] ), .S0(n3771), .S1(n3755), .Y(
        n348) );
  MXI4X1 U2736 ( .A(\regfile[12][14] ), .B(\regfile[13][14] ), .C(
        \regfile[14][14] ), .D(\regfile[15][14] ), .S0(n3772), .S1(n3742), .Y(
        n356) );
  MXI4X1 U2737 ( .A(\regfile[12][15] ), .B(\regfile[13][15] ), .C(
        \regfile[14][15] ), .D(\regfile[15][15] ), .S0(n3772), .S1(n3749), .Y(
        n364) );
  MXI4X1 U2738 ( .A(\regfile[12][16] ), .B(\regfile[13][16] ), .C(
        \regfile[14][16] ), .D(\regfile[15][16] ), .S0(n3758), .S1(n3752), .Y(
        n372) );
  MXI4X1 U2739 ( .A(\regfile[12][17] ), .B(\regfile[13][17] ), .C(
        \regfile[14][17] ), .D(\regfile[15][17] ), .S0(n3758), .S1(n3748), .Y(
        n380) );
  MXI4X1 U2740 ( .A(\regfile[12][18] ), .B(\regfile[13][18] ), .C(
        \regfile[14][18] ), .D(\regfile[15][18] ), .S0(n3759), .S1(n3742), .Y(
        n388) );
  MXI4X1 U2741 ( .A(\regfile[12][19] ), .B(\regfile[13][19] ), .C(
        \regfile[14][19] ), .D(\regfile[15][19] ), .S0(n3759), .S1(n3752), .Y(
        n396) );
  MXI4X1 U2742 ( .A(\regfile[12][20] ), .B(\regfile[13][20] ), .C(
        \regfile[14][20] ), .D(\regfile[15][20] ), .S0(n3760), .S1(n3742), .Y(
        n404) );
  MXI4X1 U2743 ( .A(\regfile[12][21] ), .B(\regfile[13][21] ), .C(
        \regfile[14][21] ), .D(\regfile[15][21] ), .S0(n3760), .S1(n3746), .Y(
        n412) );
  MXI4X1 U2744 ( .A(\regfile[12][22] ), .B(\regfile[13][22] ), .C(
        \regfile[14][22] ), .D(\regfile[15][22] ), .S0(n3761), .S1(n3744), .Y(
        n420) );
  MXI4X1 U2745 ( .A(\regfile[12][23] ), .B(\regfile[13][23] ), .C(
        \regfile[14][23] ), .D(\regfile[15][23] ), .S0(n3761), .S1(n3753), .Y(
        n428) );
  MXI4X1 U2746 ( .A(\regfile[12][24] ), .B(\regfile[13][24] ), .C(
        \regfile[14][24] ), .D(\regfile[15][24] ), .S0(n3762), .S1(n3744), .Y(
        n436) );
  MXI4X1 U2747 ( .A(\regfile[12][25] ), .B(\regfile[13][25] ), .C(
        \regfile[14][25] ), .D(\regfile[15][25] ), .S0(n3762), .S1(n3751), .Y(
        n444) );
  MXI4X1 U2748 ( .A(\regfile[12][26] ), .B(\regfile[13][26] ), .C(
        \regfile[14][26] ), .D(\regfile[15][26] ), .S0(n3763), .S1(n3751), .Y(
        n452) );
  MXI4X1 U2749 ( .A(\regfile[12][27] ), .B(\regfile[13][27] ), .C(
        \regfile[14][27] ), .D(\regfile[15][27] ), .S0(n3763), .S1(n3743), .Y(
        n460) );
  MXI4X1 U2750 ( .A(\regfile[12][28] ), .B(\regfile[13][28] ), .C(
        \regfile[14][28] ), .D(\regfile[15][28] ), .S0(n3763), .S1(n3744), .Y(
        n468) );
  MXI4X1 U2751 ( .A(\regfile[12][29] ), .B(\regfile[13][29] ), .C(
        \regfile[14][29] ), .D(\regfile[15][29] ), .S0(n3764), .S1(n3744), .Y(
        n476) );
  MXI4X1 U2752 ( .A(\regfile[12][30] ), .B(\regfile[13][30] ), .C(
        \regfile[14][30] ), .D(\regfile[15][30] ), .S0(n3764), .S1(n3744), .Y(
        n484) );
  MXI4X1 U2753 ( .A(\regfile[12][31] ), .B(\regfile[13][31] ), .C(
        \regfile[14][31] ), .D(\regfile[15][31] ), .S0(n3765), .S1(n3745), .Y(
        n492) );
  MXI4X1 U2754 ( .A(\regfile[8][0] ), .B(\regfile[9][0] ), .C(\regfile[10][0] ), .D(\regfile[11][0] ), .S0(n4290), .S1(n4278), .Y(n3846) );
  MXI4X1 U2755 ( .A(\regfile[8][1] ), .B(\regfile[9][1] ), .C(\regfile[10][1] ), .D(\regfile[11][1] ), .S0(n4291), .S1(n4275), .Y(n3854) );
  MXI4X1 U2756 ( .A(\regfile[8][2] ), .B(\regfile[9][2] ), .C(\regfile[10][2] ), .D(\regfile[11][2] ), .S0(n4291), .S1(n4268), .Y(n3862) );
  MXI4X1 U2757 ( .A(\regfile[8][3] ), .B(\regfile[9][3] ), .C(\regfile[10][3] ), .D(\regfile[11][3] ), .S0(n4292), .S1(n4271), .Y(n3870) );
  MXI4X1 U2758 ( .A(\regfile[8][4] ), .B(\regfile[9][4] ), .C(\regfile[10][4] ), .D(\regfile[11][4] ), .S0(n4292), .S1(n4271), .Y(n3878) );
  MXI4X1 U2759 ( .A(\regfile[8][5] ), .B(\regfile[9][5] ), .C(\regfile[10][5] ), .D(\regfile[11][5] ), .S0(n4293), .S1(n4271), .Y(n3886) );
  MXI4X1 U2760 ( .A(\regfile[8][6] ), .B(\regfile[9][6] ), .C(\regfile[10][6] ), .D(\regfile[11][6] ), .S0(n4293), .S1(n4272), .Y(n3894) );
  MXI4X1 U2761 ( .A(\regfile[8][7] ), .B(\regfile[9][7] ), .C(\regfile[10][7] ), .D(\regfile[11][7] ), .S0(n4294), .S1(n4272), .Y(n3902) );
  MXI4X1 U2762 ( .A(\regfile[8][8] ), .B(\regfile[9][8] ), .C(\regfile[10][8] ), .D(\regfile[11][8] ), .S0(n4294), .S1(n4272), .Y(n3910) );
  MXI4X1 U2763 ( .A(\regfile[8][9] ), .B(\regfile[9][9] ), .C(\regfile[10][9] ), .D(\regfile[11][9] ), .S0(n4295), .S1(n4273), .Y(n3918) );
  MXI4X1 U2764 ( .A(\regfile[8][10] ), .B(\regfile[9][10] ), .C(
        \regfile[10][10] ), .D(\regfile[11][10] ), .S0(n4295), .S1(n4273), .Y(
        n3926) );
  MXI4X1 U2765 ( .A(\regfile[8][11] ), .B(\regfile[9][11] ), .C(
        \regfile[10][11] ), .D(\regfile[11][11] ), .S0(n4295), .S1(n4273), .Y(
        n3934) );
  MXI4X1 U2766 ( .A(\regfile[8][12] ), .B(\regfile[9][12] ), .C(
        \regfile[10][12] ), .D(\regfile[11][12] ), .S0(n4296), .S1(n4266), .Y(
        n3942) );
  MXI4X1 U2767 ( .A(\regfile[8][13] ), .B(\regfile[9][13] ), .C(
        \regfile[10][13] ), .D(\regfile[11][13] ), .S0(n4296), .S1(n4272), .Y(
        n3950) );
  MXI4X1 U2768 ( .A(\regfile[8][14] ), .B(\regfile[9][14] ), .C(
        \regfile[10][14] ), .D(\regfile[11][14] ), .S0(n4297), .S1(n4277), .Y(
        n3958) );
  MXI4X1 U2769 ( .A(\regfile[8][15] ), .B(\regfile[9][15] ), .C(
        \regfile[10][15] ), .D(\regfile[11][15] ), .S0(n4297), .S1(n4267), .Y(
        n3966) );
  MXI4X1 U2770 ( .A(\regfile[8][16] ), .B(\regfile[9][16] ), .C(
        \regfile[10][16] ), .D(\regfile[11][16] ), .S0(n4283), .S1(n4269), .Y(
        n3974) );
  MXI4X1 U2771 ( .A(\regfile[8][17] ), .B(\regfile[9][17] ), .C(
        \regfile[10][17] ), .D(\regfile[11][17] ), .S0(n4283), .S1(n4267), .Y(
        n3982) );
  MXI4X1 U2772 ( .A(\regfile[8][18] ), .B(\regfile[9][18] ), .C(
        \regfile[10][18] ), .D(\regfile[11][18] ), .S0(n4284), .S1(n4269), .Y(
        n3990) );
  MXI4X1 U2773 ( .A(\regfile[8][19] ), .B(\regfile[9][19] ), .C(
        \regfile[10][19] ), .D(\regfile[11][19] ), .S0(n4284), .S1(n4274), .Y(
        n3998) );
  MXI4X1 U2774 ( .A(\regfile[8][20] ), .B(\regfile[9][20] ), .C(
        \regfile[10][20] ), .D(\regfile[11][20] ), .S0(n4285), .S1(n4267), .Y(
        n4006) );
  MXI4X1 U2775 ( .A(\regfile[8][21] ), .B(\regfile[9][21] ), .C(
        \regfile[10][21] ), .D(\regfile[11][21] ), .S0(n4285), .S1(n4266), .Y(
        n4014) );
  MXI4X1 U2776 ( .A(\regfile[8][22] ), .B(\regfile[9][22] ), .C(
        \regfile[10][22] ), .D(\regfile[11][22] ), .S0(n4286), .S1(n4267), .Y(
        n4022) );
  MXI4X1 U2777 ( .A(\regfile[8][23] ), .B(\regfile[9][23] ), .C(
        \regfile[10][23] ), .D(\regfile[11][23] ), .S0(n4286), .S1(n4278), .Y(
        n4030) );
  MXI4X1 U2778 ( .A(\regfile[8][24] ), .B(\regfile[9][24] ), .C(
        \regfile[10][24] ), .D(\regfile[11][24] ), .S0(n4287), .S1(n4270), .Y(
        n4038) );
  MXI4X1 U2779 ( .A(\regfile[8][25] ), .B(\regfile[9][25] ), .C(
        \regfile[10][25] ), .D(\regfile[11][25] ), .S0(n4287), .S1(n4279), .Y(
        n4046) );
  MXI4X1 U2780 ( .A(\regfile[8][26] ), .B(\regfile[9][26] ), .C(
        \regfile[10][26] ), .D(\regfile[11][26] ), .S0(n4288), .S1(n4267), .Y(
        n4054) );
  MXI4X1 U2781 ( .A(\regfile[8][27] ), .B(\regfile[9][27] ), .C(
        \regfile[10][27] ), .D(\regfile[11][27] ), .S0(n4288), .S1(n4267), .Y(
        n4062) );
  MXI4X1 U2782 ( .A(\regfile[8][28] ), .B(\regfile[9][28] ), .C(
        \regfile[10][28] ), .D(\regfile[11][28] ), .S0(n4289), .S1(n4277), .Y(
        n4070) );
  MXI4X1 U2783 ( .A(\regfile[8][29] ), .B(\regfile[9][29] ), .C(
        \regfile[10][29] ), .D(\regfile[11][29] ), .S0(n4289), .S1(n4275), .Y(
        n4078) );
  MXI4X1 U2784 ( .A(\regfile[8][30] ), .B(\regfile[9][30] ), .C(
        \regfile[10][30] ), .D(\regfile[11][30] ), .S0(n4289), .S1(n4277), .Y(
        n4086) );
  MXI4X1 U2785 ( .A(\regfile[8][31] ), .B(\regfile[9][31] ), .C(
        \regfile[10][31] ), .D(\regfile[11][31] ), .S0(n4286), .S1(n4266), .Y(
        n4094) );
  MXI4X1 U2786 ( .A(\regfile[8][0] ), .B(\regfile[9][0] ), .C(\regfile[10][0] ), .D(\regfile[11][0] ), .S0(n3765), .S1(n3745), .Y(n245) );
  MXI4X1 U2787 ( .A(\regfile[8][1] ), .B(\regfile[9][1] ), .C(\regfile[10][1] ), .D(\regfile[11][1] ), .S0(n3766), .S1(n3745), .Y(n253) );
  MXI4X1 U2788 ( .A(\regfile[8][2] ), .B(\regfile[9][2] ), .C(\regfile[10][2] ), .D(\regfile[11][2] ), .S0(n3766), .S1(n3745), .Y(n261) );
  MXI4X1 U2789 ( .A(\regfile[8][3] ), .B(\regfile[9][3] ), .C(\regfile[10][3] ), .D(\regfile[11][3] ), .S0(n3767), .S1(n3755), .Y(n269) );
  MXI4X1 U2790 ( .A(\regfile[8][4] ), .B(\regfile[9][4] ), .C(\regfile[10][4] ), .D(\regfile[11][4] ), .S0(n3767), .S1(n3753), .Y(n277) );
  MXI4X1 U2791 ( .A(\regfile[8][5] ), .B(\regfile[9][5] ), .C(\regfile[10][5] ), .D(\regfile[11][5] ), .S0(n3768), .S1(n3752), .Y(n285) );
  MXI4X1 U2792 ( .A(\regfile[8][9] ), .B(\regfile[9][9] ), .C(\regfile[10][9] ), .D(\regfile[11][9] ), .S0(n3770), .S1(n3747), .Y(n317) );
  MXI4X1 U2793 ( .A(\regfile[8][10] ), .B(\regfile[9][10] ), .C(
        \regfile[10][10] ), .D(\regfile[11][10] ), .S0(n3770), .S1(n3747), .Y(
        n325) );
  MXI4X1 U2794 ( .A(\regfile[8][11] ), .B(\regfile[9][11] ), .C(
        \regfile[10][11] ), .D(\regfile[11][11] ), .S0(n3770), .S1(n3747), .Y(
        n333) );
  MXI4X1 U2795 ( .A(\regfile[8][12] ), .B(\regfile[9][12] ), .C(
        \regfile[10][12] ), .D(\regfile[11][12] ), .S0(n3771), .S1(n3751), .Y(
        n341) );
  MXI4X1 U2796 ( .A(\regfile[8][13] ), .B(\regfile[9][13] ), .C(
        \regfile[10][13] ), .D(\regfile[11][13] ), .S0(n3771), .S1(n3742), .Y(
        n349) );
  MXI4X1 U2797 ( .A(\regfile[8][14] ), .B(\regfile[9][14] ), .C(
        \regfile[10][14] ), .D(\regfile[11][14] ), .S0(n3772), .S1(n3754), .Y(
        n357) );
  MXI4X1 U2798 ( .A(\regfile[8][15] ), .B(\regfile[9][15] ), .C(
        \regfile[10][15] ), .D(\regfile[11][15] ), .S0(n3772), .S1(n3749), .Y(
        n365) );
  MXI4X1 U2799 ( .A(\regfile[8][16] ), .B(\regfile[9][16] ), .C(
        \regfile[10][16] ), .D(\regfile[11][16] ), .S0(n3758), .S1(n3746), .Y(
        n373) );
  MXI4X1 U2800 ( .A(\regfile[8][17] ), .B(\regfile[9][17] ), .C(
        \regfile[10][17] ), .D(\regfile[11][17] ), .S0(n3758), .S1(n3743), .Y(
        n381) );
  MXI4X1 U2801 ( .A(\regfile[8][18] ), .B(\regfile[9][18] ), .C(
        \regfile[10][18] ), .D(\regfile[11][18] ), .S0(n3759), .S1(n3754), .Y(
        n389) );
  MXI4X1 U2802 ( .A(\regfile[8][19] ), .B(\regfile[9][19] ), .C(
        \regfile[10][19] ), .D(\regfile[11][19] ), .S0(n3759), .S1(n3753), .Y(
        n397) );
  MXI4X1 U2803 ( .A(\regfile[8][20] ), .B(\regfile[9][20] ), .C(
        \regfile[10][20] ), .D(\regfile[11][20] ), .S0(n3760), .S1(n3746), .Y(
        n405) );
  MXI4X1 U2804 ( .A(\regfile[8][21] ), .B(\regfile[9][21] ), .C(
        \regfile[10][21] ), .D(\regfile[11][21] ), .S0(n3760), .S1(n3752), .Y(
        n413) );
  MXI4X1 U2805 ( .A(\regfile[8][22] ), .B(\regfile[9][22] ), .C(
        \regfile[10][22] ), .D(\regfile[11][22] ), .S0(n3761), .S1(n3752), .Y(
        n421) );
  MXI4X1 U2806 ( .A(\regfile[8][23] ), .B(\regfile[9][23] ), .C(
        \regfile[10][23] ), .D(\regfile[11][23] ), .S0(n3761), .S1(n3751), .Y(
        n429) );
  MXI4X1 U2807 ( .A(\regfile[8][24] ), .B(\regfile[9][24] ), .C(
        \regfile[10][24] ), .D(\regfile[11][24] ), .S0(n3762), .S1(n3744), .Y(
        n437) );
  MXI4X1 U2808 ( .A(\regfile[8][25] ), .B(\regfile[9][25] ), .C(
        \regfile[10][25] ), .D(\regfile[11][25] ), .S0(n3762), .S1(n3752), .Y(
        n445) );
  MXI4X1 U2809 ( .A(\regfile[8][26] ), .B(\regfile[9][26] ), .C(
        \regfile[10][26] ), .D(\regfile[11][26] ), .S0(n3763), .S1(n3754), .Y(
        n453) );
  MXI4X1 U2810 ( .A(\regfile[8][27] ), .B(\regfile[9][27] ), .C(
        \regfile[10][27] ), .D(\regfile[11][27] ), .S0(n3763), .S1(n3747), .Y(
        n461) );
  MXI4X1 U2811 ( .A(\regfile[8][28] ), .B(\regfile[9][28] ), .C(
        \regfile[10][28] ), .D(\regfile[11][28] ), .S0(n3764), .S1(n3744), .Y(
        n469) );
  MXI4X1 U2812 ( .A(\regfile[8][29] ), .B(\regfile[9][29] ), .C(
        \regfile[10][29] ), .D(\regfile[11][29] ), .S0(n3764), .S1(n3744), .Y(
        n477) );
  MXI4X1 U2813 ( .A(\regfile[8][30] ), .B(\regfile[9][30] ), .C(
        \regfile[10][30] ), .D(\regfile[11][30] ), .S0(n3764), .S1(n3744), .Y(
        n485) );
  MXI4X1 U2814 ( .A(\regfile[8][31] ), .B(\regfile[9][31] ), .C(
        \regfile[10][31] ), .D(\regfile[11][31] ), .S0(n3761), .S1(n3753), .Y(
        n493) );
  NOR4X1 U2815 ( .A(Instruction[29]), .B(Instruction[28]), .C(Instruction[31]), 
        .D(Instruction[30]), .Y(n170) );
  OAI221XL U2816 ( .A0(n3657), .A1(n4367), .B0(n4952), .B1(n1793), .C0(n4577), 
        .Y(n3659) );
  OA22X1 U2817 ( .A0(n4420), .A1(n4576), .B0(n600), .B1(n4417), .Y(n4577) );
  CLKINVX1 U2818 ( .A(PCadd4[0]), .Y(n4576) );
  OAI221XL U2819 ( .A0(n3656), .A1(n4367), .B0(n4966), .B1(n1793), .C0(n4579), 
        .Y(n3660) );
  OA22X1 U2820 ( .A0(n4420), .A1(n4578), .B0(n599), .B1(n4417), .Y(n4579) );
  CLKINVX1 U2821 ( .A(PCadd4[1]), .Y(n4578) );
  OAI221XL U2822 ( .A0(n3655), .A1(n4367), .B0(n4934), .B1(n1793), .C0(n4581), 
        .Y(n3661) );
  OA22X1 U2823 ( .A0(n4420), .A1(n4580), .B0(n598), .B1(n4417), .Y(n4581) );
  OAI221XL U2824 ( .A0(n3654), .A1(n4367), .B0(n4943), .B1(n1793), .C0(n4583), 
        .Y(n3662) );
  OA22X1 U2825 ( .A0(n4420), .A1(n4582), .B0(n597), .B1(n4417), .Y(n4583) );
  OAI221XL U2826 ( .A0(n3653), .A1(n4367), .B0(n4913), .B1(n1793), .C0(n4585), 
        .Y(n3663) );
  OA22X1 U2827 ( .A0(n4420), .A1(n4584), .B0(n596), .B1(n4417), .Y(n4585) );
  OAI221XL U2828 ( .A0(n3652), .A1(n4367), .B0(n4922), .B1(n1793), .C0(n4587), 
        .Y(n3664) );
  OA22X1 U2829 ( .A0(n4420), .A1(n4586), .B0(n595), .B1(n4417), .Y(n4587) );
  CLKINVX1 U2830 ( .A(PCadd4[5]), .Y(n4586) );
  OAI221XL U2831 ( .A0(n3651), .A1(n4367), .B0(n4895), .B1(n1793), .C0(n4589), 
        .Y(n3665) );
  OA22X1 U2832 ( .A0(n4420), .A1(n4588), .B0(n594), .B1(n4417), .Y(n4589) );
  CLKINVX1 U2833 ( .A(PCadd4[6]), .Y(n4588) );
  OAI221XL U2834 ( .A0(n3650), .A1(n4367), .B0(n4904), .B1(n1793), .C0(n4591), 
        .Y(n3666) );
  OA22X1 U2835 ( .A0(n4421), .A1(n4590), .B0(n593), .B1(n4417), .Y(n4591) );
  CLKINVX1 U2836 ( .A(PCadd4[7]), .Y(n4590) );
  OAI221XL U2837 ( .A0(n3649), .A1(n4367), .B0(n4874), .B1(n1793), .C0(n4593), 
        .Y(n3667) );
  OA22X1 U2838 ( .A0(n4420), .A1(n4592), .B0(n592), .B1(n4417), .Y(n4593) );
  CLKINVX1 U2839 ( .A(PCadd4[8]), .Y(n4592) );
  OAI221XL U2840 ( .A0(n3648), .A1(n4367), .B0(n4883), .B1(n1793), .C0(n4595), 
        .Y(n3668) );
  OA22X1 U2841 ( .A0(n4420), .A1(n4594), .B0(n591), .B1(n4417), .Y(n4595) );
  CLKINVX1 U2842 ( .A(PCadd4[9]), .Y(n4594) );
  OAI221XL U2843 ( .A0(n3647), .A1(n4367), .B0(n4856), .B1(n1793), .C0(n4597), 
        .Y(n3669) );
  OA22X1 U2844 ( .A0(n4420), .A1(n4596), .B0(n590), .B1(n4417), .Y(n4597) );
  CLKINVX1 U2845 ( .A(PCadd4[10]), .Y(n4596) );
  OAI221XL U2846 ( .A0(n3646), .A1(n4367), .B0(n4865), .B1(n1793), .C0(n4599), 
        .Y(n3670) );
  OA22X1 U2847 ( .A0(n4420), .A1(n4598), .B0(n589), .B1(n4417), .Y(n4599) );
  CLKINVX1 U2848 ( .A(PCadd4[11]), .Y(n4598) );
  OAI221XL U2849 ( .A0(n3645), .A1(n4367), .B0(n4834), .B1(n1793), .C0(n4601), 
        .Y(n3671) );
  OA22X1 U2850 ( .A0(n4421), .A1(n4600), .B0(n588), .B1(n4418), .Y(n4601) );
  CLKINVX1 U2851 ( .A(PCadd4[12]), .Y(n4600) );
  OAI221XL U2852 ( .A0(n3644), .A1(n4368), .B0(n4843), .B1(n1793), .C0(n4603), 
        .Y(n3672) );
  OA22X1 U2853 ( .A0(n4421), .A1(n4602), .B0(n587), .B1(n4418), .Y(n4603) );
  CLKINVX1 U2854 ( .A(PCadd4[13]), .Y(n4602) );
  OAI221XL U2855 ( .A0(n3643), .A1(n4368), .B0(n4816), .B1(n1793), .C0(n4605), 
        .Y(n3673) );
  OA22X1 U2856 ( .A0(n4421), .A1(n4604), .B0(n586), .B1(n4418), .Y(n4605) );
  CLKINVX1 U2857 ( .A(PCadd4[14]), .Y(n4604) );
  OAI221XL U2858 ( .A0(n3642), .A1(n4368), .B0(n4825), .B1(n1793), .C0(n4607), 
        .Y(n3674) );
  OA22X1 U2859 ( .A0(n4421), .A1(n4606), .B0(n585), .B1(n4418), .Y(n4607) );
  CLKINVX1 U2860 ( .A(PCadd4[15]), .Y(n4606) );
  OAI221XL U2861 ( .A0(n3641), .A1(n4368), .B0(n4790), .B1(n1793), .C0(n4609), 
        .Y(n3675) );
  OA22X1 U2862 ( .A0(n4421), .A1(n4608), .B0(n584), .B1(n4418), .Y(n4609) );
  CLKINVX1 U2863 ( .A(PCadd4[16]), .Y(n4608) );
  OAI221XL U2864 ( .A0(n3640), .A1(n4368), .B0(n4799), .B1(n1793), .C0(n4611), 
        .Y(n3676) );
  OA22X1 U2865 ( .A0(n4421), .A1(n4610), .B0(n583), .B1(n4418), .Y(n4611) );
  CLKINVX1 U2866 ( .A(PCadd4[17]), .Y(n4610) );
  OAI221XL U2867 ( .A0(n3639), .A1(n4368), .B0(n4772), .B1(n1793), .C0(n4613), 
        .Y(n3677) );
  OA22X1 U2868 ( .A0(n4421), .A1(n4612), .B0(n582), .B1(n4418), .Y(n4613) );
  CLKINVX1 U2869 ( .A(PCadd4[18]), .Y(n4612) );
  OAI221XL U2870 ( .A0(n3638), .A1(n4368), .B0(n4781), .B1(n1793), .C0(n4615), 
        .Y(n3678) );
  OA22X1 U2871 ( .A0(n4421), .A1(n4614), .B0(n581), .B1(n4418), .Y(n4615) );
  CLKINVX1 U2872 ( .A(PCadd4[19]), .Y(n4614) );
  OAI221XL U2873 ( .A0(n3637), .A1(n4368), .B0(n4750), .B1(n1793), .C0(n4617), 
        .Y(n3679) );
  OA22X1 U2874 ( .A0(n4421), .A1(n4616), .B0(n580), .B1(n4418), .Y(n4617) );
  CLKINVX1 U2875 ( .A(PCadd4[20]), .Y(n4616) );
  OAI221XL U2876 ( .A0(n3636), .A1(n4368), .B0(n4759), .B1(n1793), .C0(n4619), 
        .Y(n3680) );
  OA22X1 U2877 ( .A0(n4421), .A1(n4618), .B0(n579), .B1(n4418), .Y(n4619) );
  CLKINVX1 U2878 ( .A(PCadd4[21]), .Y(n4618) );
  OAI221XL U2879 ( .A0(n3635), .A1(n4368), .B0(n4732), .B1(n1793), .C0(n4621), 
        .Y(n3681) );
  OA22X1 U2880 ( .A0(n4421), .A1(n4620), .B0(n578), .B1(n4418), .Y(n4621) );
  CLKINVX1 U2881 ( .A(PCadd4[22]), .Y(n4620) );
  OAI221XL U2882 ( .A0(n3634), .A1(n4368), .B0(n4741), .B1(n1793), .C0(n4623), 
        .Y(n3682) );
  OA22X1 U2883 ( .A0(n4421), .A1(n4622), .B0(n577), .B1(n4418), .Y(n4623) );
  CLKINVX1 U2884 ( .A(PCadd4[23]), .Y(n4622) );
  OAI221XL U2885 ( .A0(n3633), .A1(n4368), .B0(n4710), .B1(n1793), .C0(n4625), 
        .Y(n3683) );
  OA22X1 U2886 ( .A0(n4421), .A1(n4624), .B0(n576), .B1(n4418), .Y(n4625) );
  CLKINVX1 U2887 ( .A(PCadd4[24]), .Y(n4624) );
  OAI221XL U2888 ( .A0(n3632), .A1(n4368), .B0(n4719), .B1(n1793), .C0(n4627), 
        .Y(n3684) );
  OA22X1 U2889 ( .A0(n4421), .A1(n4626), .B0(n575), .B1(n4418), .Y(n4627) );
  CLKINVX1 U2890 ( .A(PCadd4[25]), .Y(n4626) );
  OAI221XL U2891 ( .A0(n3631), .A1(n4367), .B0(n4692), .B1(n1793), .C0(n4629), 
        .Y(n3685) );
  OA22X1 U2892 ( .A0(n4421), .A1(n4628), .B0(n574), .B1(n4418), .Y(n4629) );
  CLKINVX1 U2893 ( .A(PCadd4[26]), .Y(n4628) );
  OAI221XL U2894 ( .A0(n3630), .A1(n4368), .B0(n4701), .B1(n1793), .C0(n4631), 
        .Y(n3686) );
  OA22X1 U2895 ( .A0(n4421), .A1(n4630), .B0(n573), .B1(n4418), .Y(n4631) );
  CLKINVX1 U2896 ( .A(PCadd4[27]), .Y(n4630) );
  OAI221XL U2897 ( .A0(n3629), .A1(n4367), .B0(n4670), .B1(n1793), .C0(n4633), 
        .Y(n3687) );
  OA22X1 U2898 ( .A0(n4421), .A1(n4632), .B0(n572), .B1(n4418), .Y(n4633) );
  CLKINVX1 U2899 ( .A(PCadd4[28]), .Y(n4632) );
  OAI221XL U2900 ( .A0(n3628), .A1(n4368), .B0(n4679), .B1(n1793), .C0(n4635), 
        .Y(n3688) );
  OA22X1 U2901 ( .A0(n4421), .A1(n4634), .B0(n571), .B1(n4418), .Y(n4635) );
  CLKINVX1 U2902 ( .A(PCadd4[29]), .Y(n4634) );
  OAI221XL U2903 ( .A0(n3627), .A1(n4644), .B0(n4652), .B1(n1793), .C0(n4637), 
        .Y(n3689) );
  OA22X1 U2904 ( .A0(n4421), .A1(n4636), .B0(n570), .B1(n4418), .Y(n4637) );
  CLKINVX1 U2905 ( .A(PCadd4[30]), .Y(n4636) );
  OAI221XL U2906 ( .A0(n3626), .A1(n4644), .B0(n4661), .B1(n1793), .C0(n4642), 
        .Y(n3690) );
  OA22X1 U2907 ( .A0(n4420), .A1(n4641), .B0(n569), .B1(n4418), .Y(n4642) );
  CLKINVX1 U2908 ( .A(PCadd4[31]), .Y(n4641) );
  NOR2BX1 U2909 ( .AN(Reg_W[4]), .B(n4983), .Y(n104) );
  CLKINVX1 U2910 ( .A(n192), .Y(n4419) );
  OAI221XL U2911 ( .A0(n124), .A1(n132), .B0(n1899), .B1(MEM_RegWrite), .C0(
        n4420), .Y(n192) );
  NOR2BX2 U2912 ( .AN(Reg_W[1]), .B(Reg_W[0]), .Y(n57) );
  NOR2BX2 U2913 ( .AN(Reg_W[0]), .B(Reg_W[1]), .Y(n53) );
  NOR2X2 U2914 ( .A(Reg_W[0]), .B(Reg_W[1]), .Y(n65) );
  NOR2X1 U2915 ( .A(n4983), .B(Reg_W[4]), .Y(n61) );
  MXI2X1 U2916 ( .A(n1612), .B(n4399), .S0(n4303), .Y(n1614) );
  MXI2X1 U2917 ( .A(n1611), .B(n4410), .S0(n4303), .Y(n1616) );
  MXI2X1 U2918 ( .A(n1610), .B(n4397), .S0(n4303), .Y(n1618) );
  MXI2X1 U2919 ( .A(n1609), .B(n4398), .S0(n4303), .Y(n1620) );
  MXI2X1 U2920 ( .A(n1608), .B(n4395), .S0(n4303), .Y(n1622) );
  MXI2X1 U2921 ( .A(n1607), .B(n4396), .S0(n4303), .Y(n1624) );
  MXI2X1 U2922 ( .A(n1606), .B(n4393), .S0(n4303), .Y(n1626) );
  MXI2X1 U2923 ( .A(n1605), .B(n4394), .S0(n4303), .Y(n1628) );
  MXI2X1 U2924 ( .A(n1604), .B(n4391), .S0(n4303), .Y(n1630) );
  MXI2X1 U2925 ( .A(n1603), .B(n4392), .S0(n4303), .Y(n1632) );
  MXI2X1 U2926 ( .A(n1602), .B(n4389), .S0(n4303), .Y(n1634) );
  MXI2X1 U2927 ( .A(n1601), .B(n4390), .S0(n4303), .Y(n1636) );
  MXI2X1 U2928 ( .A(n1600), .B(n4387), .S0(n4304), .Y(n1638) );
  MXI2X1 U2929 ( .A(n1599), .B(n4388), .S0(n4304), .Y(n1640) );
  MXI2X1 U2930 ( .A(n1598), .B(n4385), .S0(n4304), .Y(n1642) );
  MXI2X1 U2931 ( .A(n1597), .B(n4386), .S0(n4304), .Y(n1644) );
  MXI2X1 U2932 ( .A(n1596), .B(n4383), .S0(n4304), .Y(n1646) );
  MXI2X1 U2933 ( .A(n1595), .B(n4384), .S0(n4304), .Y(n1648) );
  MXI2X1 U2934 ( .A(n1594), .B(n4381), .S0(n4304), .Y(n1650) );
  MXI2X1 U2935 ( .A(n1593), .B(n4382), .S0(n4304), .Y(n1652) );
  MXI2X1 U2936 ( .A(n1592), .B(n4379), .S0(n4304), .Y(n1654) );
  MXI2X1 U2937 ( .A(n1591), .B(n4380), .S0(n4304), .Y(n1656) );
  MXI2X1 U2938 ( .A(n1590), .B(n4377), .S0(n4304), .Y(n1658) );
  MXI2X1 U2939 ( .A(n1589), .B(n4378), .S0(n4304), .Y(n1660) );
  MXI2X1 U2940 ( .A(n1588), .B(n4375), .S0(n4303), .Y(n1662) );
  MXI2X1 U2941 ( .A(n1587), .B(n4376), .S0(n4304), .Y(n1664) );
  MXI2X1 U2942 ( .A(n1586), .B(n4373), .S0(n113), .Y(n1666) );
  MXI2X1 U2943 ( .A(n1585), .B(n4374), .S0(n113), .Y(n1668) );
  MXI2X1 U2944 ( .A(n1584), .B(n4371), .S0(n113), .Y(n1670) );
  MXI2X1 U2945 ( .A(n1583), .B(n4372), .S0(n113), .Y(n1672) );
  MXI2X1 U2946 ( .A(n1582), .B(n4369), .S0(n113), .Y(n1674) );
  MXI2X1 U2947 ( .A(n1581), .B(n4370), .S0(n113), .Y(n1676) );
  MXI2X1 U2948 ( .A(n1548), .B(n4399), .S0(n4307), .Y(n1742) );
  MXI2X1 U2949 ( .A(n1547), .B(n4410), .S0(n4307), .Y(n1744) );
  MXI2X1 U2950 ( .A(n1546), .B(n4397), .S0(n4307), .Y(n1746) );
  MXI2X1 U2951 ( .A(n1545), .B(n4398), .S0(n4307), .Y(n1748) );
  MXI2X1 U2952 ( .A(n1544), .B(n4395), .S0(n4307), .Y(n1750) );
  MXI2X1 U2953 ( .A(n1543), .B(n4396), .S0(n4307), .Y(n1752) );
  MXI2X1 U2954 ( .A(n1542), .B(n4393), .S0(n4307), .Y(n1754) );
  MXI2X1 U2955 ( .A(n1541), .B(n4394), .S0(n4307), .Y(n1756) );
  MXI2X1 U2956 ( .A(n1540), .B(n4391), .S0(n4307), .Y(n1758) );
  MXI2X1 U2957 ( .A(n1539), .B(n4392), .S0(n4307), .Y(n1760) );
  MXI2X1 U2958 ( .A(n1895), .B(n4389), .S0(n4307), .Y(n1762) );
  MXI2X1 U2959 ( .A(n1537), .B(n4390), .S0(n4307), .Y(n1764) );
  MXI2X1 U2960 ( .A(n1536), .B(n4387), .S0(n4308), .Y(n1766) );
  MXI2X1 U2961 ( .A(n1535), .B(n4388), .S0(n4308), .Y(n1768) );
  MXI2X1 U2962 ( .A(n1534), .B(n4385), .S0(n4308), .Y(n1770) );
  MXI2X1 U2963 ( .A(n1533), .B(n4386), .S0(n4308), .Y(n1772) );
  MXI2X1 U2964 ( .A(n1532), .B(n4383), .S0(n4308), .Y(n1774) );
  MXI2X1 U2965 ( .A(n1531), .B(n4384), .S0(n4308), .Y(n1776) );
  MXI2X1 U2966 ( .A(n1530), .B(n4381), .S0(n4308), .Y(n1778) );
  MXI2X1 U2967 ( .A(n1529), .B(n4382), .S0(n4308), .Y(n1780) );
  MXI2X1 U2968 ( .A(n1528), .B(n4379), .S0(n4308), .Y(n1782) );
  MXI2X1 U2969 ( .A(n1527), .B(n4380), .S0(n4308), .Y(n1784) );
  MXI2X1 U2970 ( .A(n1526), .B(n4377), .S0(n4308), .Y(n1786) );
  MXI2X1 U2971 ( .A(n1525), .B(n4378), .S0(n4308), .Y(n1788) );
  MXI2X1 U2972 ( .A(n1524), .B(n4375), .S0(n4307), .Y(n1790) );
  MXI2X1 U2973 ( .A(n1523), .B(n4376), .S0(n4308), .Y(n1792) );
  MXI2X1 U2974 ( .A(n1522), .B(n4373), .S0(n105), .Y(n1794) );
  MXI2X1 U2975 ( .A(n1521), .B(n4374), .S0(n105), .Y(n1796) );
  MXI2X1 U2976 ( .A(n1520), .B(n4371), .S0(n105), .Y(n1798) );
  MXI2X1 U2977 ( .A(n1519), .B(n4372), .S0(n105), .Y(n1800) );
  MXI2X1 U2978 ( .A(n1518), .B(n4369), .S0(n105), .Y(n1802) );
  MXI2X1 U2979 ( .A(n1517), .B(n4370), .S0(n105), .Y(n1804) );
  MXI2X1 U2980 ( .A(n1516), .B(n4399), .S0(n4309), .Y(n1806) );
  MXI2X1 U2981 ( .A(n1515), .B(n4410), .S0(n4309), .Y(n1808) );
  MXI2X1 U2982 ( .A(n1514), .B(n4397), .S0(n4309), .Y(n1810) );
  MXI2X1 U2983 ( .A(n1513), .B(n4398), .S0(n4309), .Y(n1812) );
  MXI2X1 U2984 ( .A(n1512), .B(n4395), .S0(n4309), .Y(n1814) );
  MXI2X1 U2985 ( .A(n1511), .B(n4396), .S0(n4309), .Y(n1816) );
  MXI2X1 U2986 ( .A(n1510), .B(n4393), .S0(n4309), .Y(n1818) );
  MXI2X1 U2987 ( .A(n1509), .B(n4394), .S0(n4309), .Y(n1820) );
  MXI2X1 U2988 ( .A(n1508), .B(n4391), .S0(n4309), .Y(n1822) );
  MXI2X1 U2989 ( .A(n1507), .B(n4392), .S0(n4309), .Y(n1824) );
  MXI2X1 U2990 ( .A(n1506), .B(n4389), .S0(n4309), .Y(n1826) );
  MXI2X1 U2991 ( .A(n1505), .B(n4390), .S0(n4309), .Y(n1828) );
  MXI2X1 U2992 ( .A(n1504), .B(n4387), .S0(n4310), .Y(n1830) );
  MXI2X1 U2993 ( .A(n1503), .B(n4388), .S0(n4310), .Y(n1832) );
  MXI2X1 U2994 ( .A(n1502), .B(n4385), .S0(n4310), .Y(n1834) );
  MXI2X1 U2995 ( .A(n1501), .B(n4386), .S0(n4310), .Y(n1836) );
  MXI2X1 U2996 ( .A(n1500), .B(n4383), .S0(n4310), .Y(n1838) );
  MXI2X1 U2997 ( .A(n1499), .B(n4384), .S0(n4310), .Y(n1840) );
  MXI2X1 U2998 ( .A(n1498), .B(n4381), .S0(n4310), .Y(n1842) );
  MXI2X1 U2999 ( .A(n1497), .B(n4382), .S0(n4310), .Y(n1844) );
  MXI2X1 U3000 ( .A(n1496), .B(n4379), .S0(n4310), .Y(n1846) );
  MXI2X1 U3001 ( .A(n1495), .B(n4380), .S0(n4310), .Y(n1848) );
  MXI2X1 U3002 ( .A(n1494), .B(n4377), .S0(n4310), .Y(n1850) );
  MXI2X1 U3003 ( .A(n1493), .B(n4378), .S0(n4310), .Y(n1852) );
  MXI2X1 U3004 ( .A(n1492), .B(n4375), .S0(n4309), .Y(n1854) );
  MXI2X1 U3005 ( .A(n1491), .B(n4376), .S0(n4310), .Y(n1856) );
  MXI2X1 U3006 ( .A(n1490), .B(n4373), .S0(n115), .Y(n1858) );
  MXI2X1 U3007 ( .A(n1489), .B(n4374), .S0(n115), .Y(n1860) );
  MXI2X1 U3008 ( .A(n1488), .B(n4371), .S0(n115), .Y(n1862) );
  MXI2X1 U3009 ( .A(n1487), .B(n4372), .S0(n115), .Y(n1864) );
  MXI2X1 U3010 ( .A(n1486), .B(n4369), .S0(n115), .Y(n1866) );
  MXI2X1 U3011 ( .A(n1485), .B(n4370), .S0(n115), .Y(n1868) );
  MXI2X1 U3012 ( .A(n1484), .B(n4399), .S0(n4311), .Y(n1870) );
  MXI2X1 U3013 ( .A(n1483), .B(n4410), .S0(n4311), .Y(n1872) );
  MXI2X1 U3014 ( .A(n1482), .B(n4397), .S0(n4311), .Y(n1874) );
  MXI2X1 U3015 ( .A(n1481), .B(n4398), .S0(n4311), .Y(n1876) );
  MXI2X1 U3016 ( .A(n1480), .B(n4395), .S0(n4311), .Y(n1878) );
  MXI2X1 U3017 ( .A(n1479), .B(n4396), .S0(n4311), .Y(n1880) );
  MXI2X1 U3018 ( .A(n1478), .B(n4393), .S0(n4311), .Y(n1882) );
  MXI2X1 U3019 ( .A(n1477), .B(n4394), .S0(n4311), .Y(n1884) );
  MXI2X1 U3020 ( .A(n1476), .B(n4391), .S0(n4311), .Y(n1886) );
  MXI2X1 U3021 ( .A(n1475), .B(n4392), .S0(n4311), .Y(n1888) );
  MXI2X1 U3022 ( .A(n1474), .B(n4389), .S0(n4311), .Y(n1890) );
  MXI2X1 U3023 ( .A(n1473), .B(n4390), .S0(n4311), .Y(n1892) );
  MXI2X1 U3024 ( .A(n1472), .B(n4387), .S0(n4312), .Y(n1894) );
  MXI2X1 U3025 ( .A(n1471), .B(n4388), .S0(n4312), .Y(n1896) );
  MXI2X1 U3026 ( .A(n1470), .B(n4385), .S0(n4312), .Y(n1898) );
  MXI2X1 U3027 ( .A(n1469), .B(n4386), .S0(n4312), .Y(n1900) );
  MXI2X1 U3028 ( .A(n1468), .B(n4383), .S0(n4312), .Y(n1902) );
  MXI2X1 U3029 ( .A(n1467), .B(n4384), .S0(n4312), .Y(n1904) );
  MXI2X1 U3030 ( .A(n1466), .B(n4381), .S0(n4312), .Y(n1906) );
  MXI2X1 U3031 ( .A(n1465), .B(n4382), .S0(n4312), .Y(n1908) );
  MXI2X1 U3032 ( .A(n1464), .B(n4379), .S0(n4312), .Y(n1910) );
  MXI2X1 U3033 ( .A(n1463), .B(n4380), .S0(n4312), .Y(n1912) );
  MXI2X1 U3034 ( .A(n1462), .B(n4377), .S0(n4312), .Y(n1914) );
  MXI2X1 U3035 ( .A(n1461), .B(n4378), .S0(n4312), .Y(n1916) );
  MXI2X1 U3036 ( .A(n1460), .B(n4375), .S0(n4311), .Y(n1918) );
  MXI2X1 U3037 ( .A(n1459), .B(n4376), .S0(n4312), .Y(n1920) );
  MXI2X1 U3038 ( .A(n1458), .B(n4373), .S0(n135), .Y(n1922) );
  MXI2X1 U3039 ( .A(n1457), .B(n4374), .S0(n135), .Y(n1924) );
  MXI2X1 U3040 ( .A(n1456), .B(n4371), .S0(n135), .Y(n1926) );
  MXI2X1 U3041 ( .A(n1455), .B(n4372), .S0(n135), .Y(n1928) );
  MXI2X1 U3042 ( .A(n1454), .B(n4369), .S0(n135), .Y(n1930) );
  MXI2X1 U3043 ( .A(n1453), .B(n4370), .S0(n135), .Y(n1932) );
  MXI2X1 U3044 ( .A(n1452), .B(n4399), .S0(n4313), .Y(n1934) );
  MXI2X1 U3045 ( .A(n1451), .B(n4410), .S0(n4313), .Y(n1936) );
  MXI2X1 U3046 ( .A(n1450), .B(n4397), .S0(n4313), .Y(n1938) );
  MXI2X1 U3047 ( .A(n1449), .B(n4398), .S0(n4313), .Y(n1940) );
  MXI2X1 U3048 ( .A(n1448), .B(n4395), .S0(n4313), .Y(n1942) );
  MXI2X1 U3049 ( .A(n1447), .B(n4396), .S0(n4313), .Y(n1944) );
  MXI2X1 U3050 ( .A(n1446), .B(n4393), .S0(n4313), .Y(n1946) );
  MXI2X1 U3051 ( .A(n1445), .B(n4394), .S0(n4313), .Y(n1948) );
  MXI2X1 U3052 ( .A(n1444), .B(n4391), .S0(n4313), .Y(n1950) );
  MXI2X1 U3053 ( .A(n1443), .B(n4392), .S0(n4313), .Y(n1952) );
  MXI2X1 U3054 ( .A(n1442), .B(n4389), .S0(n4313), .Y(n1954) );
  MXI2X1 U3055 ( .A(n1441), .B(n4390), .S0(n4313), .Y(n1956) );
  MXI2X1 U3056 ( .A(n1440), .B(n4387), .S0(n4314), .Y(n1958) );
  MXI2X1 U3057 ( .A(n1439), .B(n4388), .S0(n4314), .Y(n1960) );
  MXI2X1 U3058 ( .A(n1438), .B(n4385), .S0(n4314), .Y(n1962) );
  MXI2X1 U3059 ( .A(n1437), .B(n4386), .S0(n4314), .Y(n1964) );
  MXI2X1 U3060 ( .A(n1436), .B(n4383), .S0(n4314), .Y(n1966) );
  MXI2X1 U3061 ( .A(n1435), .B(n4384), .S0(n4314), .Y(n1968) );
  MXI2X1 U3062 ( .A(n1434), .B(n4381), .S0(n4314), .Y(n1970) );
  MXI2X1 U3063 ( .A(n1433), .B(n4382), .S0(n4314), .Y(n1972) );
  MXI2X1 U3064 ( .A(n1432), .B(n4379), .S0(n4314), .Y(n1974) );
  MXI2X1 U3065 ( .A(n1431), .B(n4380), .S0(n4314), .Y(n1976) );
  MXI2X1 U3066 ( .A(n1430), .B(n4377), .S0(n4314), .Y(n1978) );
  MXI2X1 U3067 ( .A(n1429), .B(n4378), .S0(n4314), .Y(n1980) );
  MXI2X1 U3068 ( .A(n1428), .B(n4375), .S0(n4313), .Y(n1982) );
  MXI2X1 U3069 ( .A(n1427), .B(n4376), .S0(n4314), .Y(n1984) );
  MXI2X1 U3070 ( .A(n1426), .B(n4373), .S0(n126), .Y(n1986) );
  MXI2X1 U3071 ( .A(n1425), .B(n4374), .S0(n126), .Y(n1988) );
  MXI2X1 U3072 ( .A(n1424), .B(n4371), .S0(n126), .Y(n1990) );
  MXI2X1 U3073 ( .A(n1423), .B(n4372), .S0(n126), .Y(n1992) );
  MXI2X1 U3074 ( .A(n1422), .B(n4369), .S0(n126), .Y(n1994) );
  MXI2X1 U3075 ( .A(n1421), .B(n4370), .S0(n126), .Y(n1996) );
  MXI2X1 U3076 ( .A(n1420), .B(n4399), .S0(n4315), .Y(n1998) );
  MXI2X1 U3077 ( .A(n1419), .B(n4410), .S0(n4315), .Y(n2000) );
  MXI2X1 U3078 ( .A(n1418), .B(n4397), .S0(n4315), .Y(n2002) );
  MXI2X1 U3079 ( .A(n1417), .B(n4398), .S0(n4315), .Y(n2004) );
  MXI2X1 U3080 ( .A(n1416), .B(n4395), .S0(n4315), .Y(n2006) );
  MXI2X1 U3081 ( .A(n1415), .B(n4396), .S0(n4315), .Y(n2008) );
  MXI2X1 U3082 ( .A(n1414), .B(n4393), .S0(n4315), .Y(n2010) );
  MXI2X1 U3083 ( .A(n1413), .B(n4394), .S0(n4315), .Y(n2012) );
  MXI2X1 U3084 ( .A(n1412), .B(n4391), .S0(n4315), .Y(n2014) );
  MXI2X1 U3085 ( .A(n1411), .B(n4392), .S0(n4315), .Y(n2016) );
  MXI2X1 U3086 ( .A(n1410), .B(n4389), .S0(n4315), .Y(n2018) );
  MXI2X1 U3087 ( .A(n1409), .B(n4390), .S0(n4315), .Y(n2020) );
  MXI2X1 U3088 ( .A(n1408), .B(n4387), .S0(n4316), .Y(n2022) );
  MXI2X1 U3089 ( .A(n1407), .B(n4388), .S0(n4316), .Y(n2024) );
  MXI2X1 U3090 ( .A(n1406), .B(n4385), .S0(n4316), .Y(n2026) );
  MXI2X1 U3091 ( .A(n1405), .B(n4386), .S0(n4316), .Y(n2028) );
  MXI2X1 U3092 ( .A(n1404), .B(n4383), .S0(n4316), .Y(n2030) );
  MXI2X1 U3093 ( .A(n1403), .B(n4384), .S0(n4316), .Y(n2032) );
  MXI2X1 U3094 ( .A(n1402), .B(n4381), .S0(n4316), .Y(n2034) );
  MXI2X1 U3095 ( .A(n1401), .B(n4382), .S0(n4316), .Y(n2036) );
  MXI2X1 U3096 ( .A(n1400), .B(n4379), .S0(n4316), .Y(n2038) );
  MXI2X1 U3097 ( .A(n1399), .B(n4380), .S0(n4316), .Y(n2040) );
  MXI2X1 U3098 ( .A(n1398), .B(n4377), .S0(n4316), .Y(n2042) );
  MXI2X1 U3099 ( .A(n1397), .B(n4378), .S0(n4316), .Y(n2044) );
  MXI2X1 U3100 ( .A(n1396), .B(n4375), .S0(n4315), .Y(n2046) );
  MXI2X1 U3101 ( .A(n1395), .B(n4376), .S0(n4316), .Y(n2048) );
  MXI2X1 U3102 ( .A(n1394), .B(n4373), .S0(n106), .Y(n2050) );
  MXI2X1 U3103 ( .A(n1393), .B(n4374), .S0(n106), .Y(n2052) );
  MXI2X1 U3104 ( .A(n1392), .B(n4371), .S0(n106), .Y(n2054) );
  MXI2X1 U3105 ( .A(n1391), .B(n4372), .S0(n106), .Y(n2056) );
  MXI2X1 U3106 ( .A(n1390), .B(n4369), .S0(n106), .Y(n2058) );
  MXI2X1 U3107 ( .A(n1389), .B(n4370), .S0(n106), .Y(n2060) );
  MXI2X1 U3108 ( .A(n1388), .B(n4399), .S0(n4317), .Y(n2062) );
  MXI2X1 U3109 ( .A(n1387), .B(n4410), .S0(n4317), .Y(n2064) );
  MXI2X1 U3110 ( .A(n1386), .B(n4397), .S0(n4317), .Y(n2066) );
  MXI2X1 U3111 ( .A(n1385), .B(n4398), .S0(n4317), .Y(n2068) );
  MXI2X1 U3112 ( .A(n1384), .B(n4395), .S0(n4317), .Y(n2070) );
  MXI2X1 U3113 ( .A(n1383), .B(n4396), .S0(n4317), .Y(n2072) );
  MXI2X1 U3114 ( .A(n1382), .B(n4393), .S0(n4317), .Y(n2074) );
  MXI2X1 U3115 ( .A(n1381), .B(n4394), .S0(n4317), .Y(n2076) );
  MXI2X1 U3116 ( .A(n1380), .B(n4391), .S0(n4317), .Y(n2078) );
  MXI2X1 U3117 ( .A(n1379), .B(n4392), .S0(n4317), .Y(n2080) );
  MXI2X1 U3118 ( .A(n1378), .B(n4389), .S0(n4317), .Y(n2082) );
  MXI2X1 U3119 ( .A(n1377), .B(n4390), .S0(n4317), .Y(n2084) );
  MXI2X1 U3120 ( .A(n1376), .B(n4387), .S0(n4318), .Y(n2086) );
  MXI2X1 U3121 ( .A(n1375), .B(n4388), .S0(n4318), .Y(n2088) );
  MXI2X1 U3122 ( .A(n1374), .B(n4385), .S0(n4318), .Y(n2090) );
  MXI2X1 U3123 ( .A(n1373), .B(n4386), .S0(n4318), .Y(n2092) );
  MXI2X1 U3124 ( .A(n1372), .B(n4383), .S0(n4318), .Y(n2094) );
  MXI2X1 U3125 ( .A(n1371), .B(n4384), .S0(n4318), .Y(n2096) );
  MXI2X1 U3126 ( .A(n1370), .B(n4381), .S0(n4318), .Y(n2098) );
  MXI2X1 U3127 ( .A(n1369), .B(n4382), .S0(n4318), .Y(n2100) );
  MXI2X1 U3128 ( .A(n1368), .B(n4379), .S0(n4318), .Y(n2102) );
  MXI2X1 U3129 ( .A(n1367), .B(n4380), .S0(n4318), .Y(n2104) );
  MXI2X1 U3130 ( .A(n1366), .B(n4377), .S0(n4318), .Y(n2106) );
  MXI2X1 U3131 ( .A(n1365), .B(n4378), .S0(n4318), .Y(n2108) );
  MXI2X1 U3132 ( .A(n1364), .B(n4375), .S0(n4317), .Y(n2110) );
  MXI2X1 U3133 ( .A(n1363), .B(n4376), .S0(n4318), .Y(n2112) );
  MXI2X1 U3134 ( .A(n1362), .B(n4373), .S0(n116), .Y(n2114) );
  MXI2X1 U3135 ( .A(n1361), .B(n4374), .S0(n116), .Y(n2116) );
  MXI2X1 U3136 ( .A(n1360), .B(n4371), .S0(n116), .Y(n2118) );
  MXI2X1 U3137 ( .A(n1359), .B(n4372), .S0(n116), .Y(n2120) );
  MXI2X1 U3138 ( .A(n1358), .B(n4369), .S0(n116), .Y(n2122) );
  MXI2X1 U3139 ( .A(n1357), .B(n4370), .S0(n116), .Y(n2124) );
  MXI2X1 U3140 ( .A(n1356), .B(n4399), .S0(n4319), .Y(n2126) );
  MXI2X1 U3141 ( .A(n1355), .B(n4410), .S0(n4319), .Y(n2128) );
  MXI2X1 U3142 ( .A(n1354), .B(n4397), .S0(n4319), .Y(n2130) );
  MXI2X1 U3143 ( .A(n1353), .B(n4398), .S0(n4319), .Y(n2132) );
  MXI2X1 U3144 ( .A(n1352), .B(n4395), .S0(n4319), .Y(n2134) );
  MXI2X1 U3145 ( .A(n1351), .B(n4396), .S0(n4319), .Y(n2136) );
  MXI2X1 U3146 ( .A(n1350), .B(n4393), .S0(n4319), .Y(n2138) );
  MXI2X1 U3147 ( .A(n1349), .B(n4394), .S0(n4319), .Y(n2140) );
  MXI2X1 U3148 ( .A(n1348), .B(n4391), .S0(n4319), .Y(n2142) );
  MXI2X1 U3149 ( .A(n1347), .B(n4392), .S0(n4319), .Y(n2144) );
  MXI2X1 U3150 ( .A(n1346), .B(n4389), .S0(n4319), .Y(n2146) );
  MXI2X1 U3151 ( .A(n1345), .B(n4390), .S0(n4319), .Y(n2148) );
  MXI2X1 U3152 ( .A(n1344), .B(n4387), .S0(n4320), .Y(n2150) );
  MXI2X1 U3153 ( .A(n1343), .B(n4388), .S0(n4320), .Y(n2152) );
  MXI2X1 U3154 ( .A(n1342), .B(n4385), .S0(n4320), .Y(n2154) );
  MXI2X1 U3155 ( .A(n1341), .B(n4386), .S0(n4320), .Y(n2156) );
  MXI2X1 U3156 ( .A(n1340), .B(n4383), .S0(n4320), .Y(n2158) );
  MXI2X1 U3157 ( .A(n1339), .B(n4384), .S0(n4320), .Y(n2160) );
  MXI2X1 U3158 ( .A(n1338), .B(n4381), .S0(n4320), .Y(n2162) );
  MXI2X1 U3159 ( .A(n1337), .B(n4382), .S0(n4320), .Y(n2164) );
  MXI2X1 U3160 ( .A(n1336), .B(n4379), .S0(n4320), .Y(n2166) );
  MXI2X1 U3161 ( .A(n1335), .B(n4380), .S0(n4320), .Y(n2168) );
  MXI2X1 U3162 ( .A(n1334), .B(n4377), .S0(n4320), .Y(n2170) );
  MXI2X1 U3163 ( .A(n1333), .B(n4378), .S0(n4320), .Y(n2172) );
  MXI2X1 U3164 ( .A(n1332), .B(n4375), .S0(n4319), .Y(n2174) );
  MXI2X1 U3165 ( .A(n1331), .B(n4376), .S0(n4320), .Y(n2176) );
  MXI2X1 U3166 ( .A(n1330), .B(n4373), .S0(n136), .Y(n2178) );
  MXI2X1 U3167 ( .A(n1329), .B(n4374), .S0(n136), .Y(n2180) );
  MXI2X1 U3168 ( .A(n1328), .B(n4371), .S0(n136), .Y(n2182) );
  MXI2X1 U3169 ( .A(n1327), .B(n4372), .S0(n136), .Y(n2184) );
  MXI2X1 U3170 ( .A(n1326), .B(n4369), .S0(n136), .Y(n2186) );
  MXI2X1 U3171 ( .A(n1325), .B(n4370), .S0(n136), .Y(n2188) );
  MXI2X1 U3172 ( .A(n1324), .B(n4399), .S0(n4321), .Y(n2190) );
  MXI2X1 U3173 ( .A(n1323), .B(n4410), .S0(n4321), .Y(n2192) );
  MXI2X1 U3174 ( .A(n1322), .B(n4397), .S0(n4321), .Y(n2194) );
  MXI2X1 U3175 ( .A(n1321), .B(n4398), .S0(n4321), .Y(n2196) );
  MXI2X1 U3176 ( .A(n1320), .B(n4395), .S0(n4321), .Y(n2198) );
  MXI2X1 U3177 ( .A(n1319), .B(n4396), .S0(n4321), .Y(n2200) );
  MXI2X1 U3178 ( .A(n1318), .B(n4393), .S0(n4321), .Y(n2202) );
  MXI2X1 U3179 ( .A(n1317), .B(n4394), .S0(n4321), .Y(n2204) );
  MXI2X1 U3180 ( .A(n1316), .B(n4391), .S0(n4321), .Y(n2206) );
  MXI2X1 U3181 ( .A(n1315), .B(n4392), .S0(n4321), .Y(n2208) );
  MXI2X1 U3182 ( .A(n1314), .B(n4389), .S0(n4321), .Y(n2210) );
  MXI2X1 U3183 ( .A(n1313), .B(n4390), .S0(n4321), .Y(n2212) );
  MXI2X1 U3184 ( .A(n1312), .B(n4387), .S0(n4322), .Y(n2214) );
  MXI2X1 U3185 ( .A(n1311), .B(n4388), .S0(n4322), .Y(n2216) );
  MXI2X1 U3186 ( .A(n1310), .B(n4385), .S0(n4322), .Y(n2218) );
  MXI2X1 U3187 ( .A(n1309), .B(n4386), .S0(n4322), .Y(n2220) );
  MXI2X1 U3188 ( .A(n1308), .B(n4383), .S0(n4322), .Y(n2222) );
  MXI2X1 U3189 ( .A(n1307), .B(n4384), .S0(n4322), .Y(n2224) );
  MXI2X1 U3190 ( .A(n1306), .B(n4381), .S0(n4322), .Y(n2226) );
  MXI2X1 U3191 ( .A(n1305), .B(n4382), .S0(n4322), .Y(n2228) );
  MXI2X1 U3192 ( .A(n1304), .B(n4379), .S0(n4322), .Y(n2230) );
  MXI2X1 U3193 ( .A(n1303), .B(n4380), .S0(n4322), .Y(n2232) );
  MXI2X1 U3194 ( .A(n1302), .B(n4377), .S0(n4322), .Y(n2234) );
  MXI2X1 U3195 ( .A(n1301), .B(n4378), .S0(n4322), .Y(n2236) );
  MXI2X1 U3196 ( .A(n1300), .B(n4375), .S0(n4321), .Y(n2238) );
  MXI2X1 U3197 ( .A(n1299), .B(n4376), .S0(n4322), .Y(n2240) );
  MXI2X1 U3198 ( .A(n1298), .B(n4373), .S0(n127), .Y(n2242) );
  MXI2X1 U3199 ( .A(n1297), .B(n4374), .S0(n127), .Y(n2244) );
  MXI2X1 U3200 ( .A(n1296), .B(n4371), .S0(n127), .Y(n2246) );
  MXI2X1 U3201 ( .A(n1295), .B(n4372), .S0(n127), .Y(n2248) );
  MXI2X1 U3202 ( .A(n1294), .B(n4369), .S0(n127), .Y(n2250) );
  MXI2X1 U3203 ( .A(n1293), .B(n4370), .S0(n127), .Y(n2252) );
  MXI2X1 U3204 ( .A(n1292), .B(n4399), .S0(n4323), .Y(n2254) );
  MXI2X1 U3205 ( .A(n1291), .B(n4410), .S0(n4323), .Y(n2256) );
  MXI2X1 U3206 ( .A(n1290), .B(n4397), .S0(n4323), .Y(n2258) );
  MXI2X1 U3207 ( .A(n1289), .B(n4398), .S0(n4323), .Y(n2260) );
  MXI2X1 U3208 ( .A(n1288), .B(n4395), .S0(n4323), .Y(n2262) );
  MXI2X1 U3209 ( .A(n1287), .B(n4396), .S0(n4323), .Y(n2264) );
  MXI2X1 U3210 ( .A(n1286), .B(n4393), .S0(n4323), .Y(n2266) );
  MXI2X1 U3211 ( .A(n1285), .B(n4394), .S0(n4323), .Y(n2268) );
  MXI2X1 U3212 ( .A(n1284), .B(n4391), .S0(n4323), .Y(n2270) );
  MXI2X1 U3213 ( .A(n1283), .B(n4392), .S0(n4323), .Y(n2272) );
  MXI2X1 U3214 ( .A(n1282), .B(n4389), .S0(n4323), .Y(n2274) );
  MXI2X1 U3215 ( .A(n1281), .B(n4390), .S0(n4323), .Y(n2276) );
  MXI2X1 U3216 ( .A(n1280), .B(n4387), .S0(n4324), .Y(n2278) );
  MXI2X1 U3217 ( .A(n1279), .B(n4388), .S0(n4324), .Y(n2280) );
  MXI2X1 U3218 ( .A(n1278), .B(n4385), .S0(n4324), .Y(n2282) );
  MXI2X1 U3219 ( .A(n1277), .B(n4386), .S0(n4324), .Y(n2284) );
  MXI2X1 U3220 ( .A(n1276), .B(n4383), .S0(n4324), .Y(n2286) );
  MXI2X1 U3221 ( .A(n1275), .B(n4384), .S0(n4324), .Y(n2288) );
  MXI2X1 U3222 ( .A(n1274), .B(n4381), .S0(n4324), .Y(n2290) );
  MXI2X1 U3223 ( .A(n1273), .B(n4382), .S0(n4324), .Y(n2292) );
  MXI2X1 U3224 ( .A(n1272), .B(n4379), .S0(n4324), .Y(n2294) );
  MXI2X1 U3225 ( .A(n1271), .B(n4380), .S0(n4324), .Y(n2296) );
  MXI2X1 U3226 ( .A(n1270), .B(n4377), .S0(n4324), .Y(n2298) );
  MXI2X1 U3227 ( .A(n1269), .B(n4378), .S0(n4324), .Y(n2300) );
  MXI2X1 U3228 ( .A(n1268), .B(n4375), .S0(n4323), .Y(n2302) );
  MXI2X1 U3229 ( .A(n1267), .B(n4376), .S0(n4324), .Y(n2304) );
  MXI2X1 U3230 ( .A(n1266), .B(n4373), .S0(n108), .Y(n2306) );
  MXI2X1 U3231 ( .A(n1265), .B(n4374), .S0(n108), .Y(n2308) );
  MXI2X1 U3232 ( .A(n1264), .B(n4371), .S0(n108), .Y(n2310) );
  MXI2X1 U3233 ( .A(n1263), .B(n4372), .S0(n108), .Y(n2312) );
  MXI2X1 U3234 ( .A(n1262), .B(n4369), .S0(n108), .Y(n2314) );
  MXI2X1 U3235 ( .A(n1261), .B(n4370), .S0(n108), .Y(n2316) );
  MXI2X1 U3236 ( .A(n1260), .B(n4399), .S0(n4325), .Y(n2318) );
  MXI2X1 U3237 ( .A(n1259), .B(n4410), .S0(n4325), .Y(n2320) );
  MXI2X1 U3238 ( .A(n1258), .B(n4397), .S0(n4325), .Y(n2322) );
  MXI2X1 U3239 ( .A(n1257), .B(n4398), .S0(n4325), .Y(n2324) );
  MXI2X1 U3240 ( .A(n1256), .B(n4395), .S0(n4325), .Y(n2326) );
  MXI2X1 U3241 ( .A(n1255), .B(n4396), .S0(n4325), .Y(n2328) );
  MXI2X1 U3242 ( .A(n1254), .B(n4393), .S0(n4325), .Y(n2330) );
  MXI2X1 U3243 ( .A(n1253), .B(n4394), .S0(n4325), .Y(n2332) );
  MXI2X1 U3244 ( .A(n1252), .B(n4391), .S0(n4325), .Y(n2334) );
  MXI2X1 U3245 ( .A(n1251), .B(n4392), .S0(n4325), .Y(n2336) );
  MXI2X1 U3246 ( .A(n1250), .B(n4389), .S0(n4325), .Y(n2338) );
  MXI2X1 U3247 ( .A(n1249), .B(n4390), .S0(n4325), .Y(n2340) );
  MXI2X1 U3248 ( .A(n1248), .B(n4387), .S0(n4326), .Y(n2342) );
  MXI2X1 U3249 ( .A(n1247), .B(n4388), .S0(n4326), .Y(n2344) );
  MXI2X1 U3250 ( .A(n1246), .B(n4385), .S0(n4326), .Y(n2346) );
  MXI2X1 U3251 ( .A(n1245), .B(n4386), .S0(n4326), .Y(n2348) );
  MXI2X1 U3252 ( .A(n1244), .B(n4383), .S0(n4326), .Y(n2350) );
  MXI2X1 U3253 ( .A(n1243), .B(n4384), .S0(n4326), .Y(n2352) );
  MXI2X1 U3254 ( .A(n1242), .B(n4381), .S0(n4326), .Y(n2354) );
  MXI2X1 U3255 ( .A(n1241), .B(n4382), .S0(n4326), .Y(n2356) );
  MXI2X1 U3256 ( .A(n1240), .B(n4379), .S0(n4326), .Y(n2358) );
  MXI2X1 U3257 ( .A(n1239), .B(n4380), .S0(n4326), .Y(n2360) );
  MXI2X1 U3258 ( .A(n1238), .B(n4377), .S0(n4326), .Y(n2362) );
  MXI2X1 U3259 ( .A(n1237), .B(n4378), .S0(n4326), .Y(n2364) );
  MXI2X1 U3260 ( .A(n1236), .B(n4375), .S0(n4325), .Y(n2366) );
  MXI2X1 U3261 ( .A(n1235), .B(n4376), .S0(n4326), .Y(n2368) );
  MXI2X1 U3262 ( .A(n1234), .B(n4373), .S0(n118), .Y(n2370) );
  MXI2X1 U3263 ( .A(n1233), .B(n4374), .S0(n118), .Y(n2372) );
  MXI2X1 U3264 ( .A(n1232), .B(n4371), .S0(n118), .Y(n2374) );
  MXI2X1 U3265 ( .A(n1231), .B(n4372), .S0(n118), .Y(n2376) );
  MXI2X1 U3266 ( .A(n1230), .B(n4369), .S0(n118), .Y(n2378) );
  MXI2X1 U3267 ( .A(n1229), .B(n4370), .S0(n118), .Y(n2380) );
  MXI2X1 U3268 ( .A(n1228), .B(n4399), .S0(n4327), .Y(n2382) );
  MXI2X1 U3269 ( .A(n1227), .B(n4410), .S0(n4327), .Y(n2384) );
  MXI2X1 U3270 ( .A(n1226), .B(n4397), .S0(n4327), .Y(n2386) );
  MXI2X1 U3271 ( .A(n1225), .B(n4398), .S0(n4327), .Y(n2388) );
  MXI2X1 U3272 ( .A(n1224), .B(n4395), .S0(n4327), .Y(n2390) );
  MXI2X1 U3273 ( .A(n1223), .B(n4396), .S0(n4327), .Y(n2392) );
  MXI2X1 U3274 ( .A(n1222), .B(n4393), .S0(n4327), .Y(n2394) );
  MXI2X1 U3275 ( .A(n1221), .B(n4394), .S0(n4327), .Y(n2396) );
  MXI2X1 U3276 ( .A(n1220), .B(n4391), .S0(n4327), .Y(n2398) );
  MXI2X1 U3277 ( .A(n1219), .B(n4392), .S0(n4327), .Y(n2400) );
  MXI2X1 U3278 ( .A(n1218), .B(n4389), .S0(n4327), .Y(n2402) );
  MXI2X1 U3279 ( .A(n1217), .B(n4390), .S0(n4327), .Y(n2404) );
  MXI2X1 U3280 ( .A(n1216), .B(n4387), .S0(n4328), .Y(n2406) );
  MXI2X1 U3281 ( .A(n1215), .B(n4388), .S0(n4328), .Y(n2408) );
  MXI2X1 U3282 ( .A(n1214), .B(n4385), .S0(n4328), .Y(n2410) );
  MXI2X1 U3283 ( .A(n1213), .B(n4386), .S0(n4328), .Y(n2412) );
  MXI2X1 U3284 ( .A(n1212), .B(n4383), .S0(n4328), .Y(n2414) );
  MXI2X1 U3285 ( .A(n1211), .B(n4384), .S0(n4328), .Y(n2416) );
  MXI2X1 U3286 ( .A(n1210), .B(n4381), .S0(n4328), .Y(n2418) );
  MXI2X1 U3287 ( .A(n1209), .B(n4382), .S0(n4328), .Y(n2420) );
  MXI2X1 U3288 ( .A(n1208), .B(n4379), .S0(n4328), .Y(n2422) );
  MXI2X1 U3289 ( .A(n1207), .B(n4380), .S0(n4328), .Y(n2424) );
  MXI2X1 U3290 ( .A(n1206), .B(n4377), .S0(n4328), .Y(n2426) );
  MXI2X1 U3291 ( .A(n1205), .B(n4378), .S0(n4328), .Y(n2428) );
  MXI2X1 U3292 ( .A(n1204), .B(n4375), .S0(n4327), .Y(n2430) );
  MXI2X1 U3293 ( .A(n1203), .B(n4376), .S0(n4328), .Y(n2432) );
  MXI2X1 U3294 ( .A(n1202), .B(n4373), .S0(n137), .Y(n2434) );
  MXI2X1 U3295 ( .A(n1201), .B(n4374), .S0(n137), .Y(n2436) );
  MXI2X1 U3296 ( .A(n1200), .B(n4371), .S0(n137), .Y(n2438) );
  MXI2X1 U3297 ( .A(n1199), .B(n4372), .S0(n137), .Y(n2440) );
  MXI2X1 U3298 ( .A(n1198), .B(n4369), .S0(n137), .Y(n2442) );
  MXI2X1 U3299 ( .A(n1197), .B(n4370), .S0(n137), .Y(n2444) );
  MXI2X1 U3300 ( .A(n1196), .B(n4399), .S0(n4329), .Y(n2446) );
  MXI2X1 U3301 ( .A(n1195), .B(n4410), .S0(n4329), .Y(n2448) );
  MXI2X1 U3302 ( .A(n1194), .B(n4397), .S0(n4329), .Y(n2450) );
  MXI2X1 U3303 ( .A(n1193), .B(n4398), .S0(n4329), .Y(n2452) );
  MXI2X1 U3304 ( .A(n1192), .B(n4395), .S0(n4329), .Y(n2454) );
  MXI2X1 U3305 ( .A(n1191), .B(n4396), .S0(n4329), .Y(n2456) );
  MXI2X1 U3306 ( .A(n1190), .B(n4393), .S0(n4329), .Y(n2458) );
  MXI2X1 U3307 ( .A(n1189), .B(n4394), .S0(n4329), .Y(n2460) );
  MXI2X1 U3308 ( .A(n1188), .B(n4391), .S0(n4329), .Y(n2462) );
  MXI2X1 U3309 ( .A(n1187), .B(n4392), .S0(n4329), .Y(n2464) );
  MXI2X1 U3310 ( .A(n1186), .B(n4389), .S0(n4329), .Y(n2466) );
  MXI2X1 U3311 ( .A(n1185), .B(n4390), .S0(n4329), .Y(n2468) );
  MXI2X1 U3312 ( .A(n1184), .B(n4387), .S0(n4330), .Y(n2470) );
  MXI2X1 U3313 ( .A(n1183), .B(n4388), .S0(n4330), .Y(n2472) );
  MXI2X1 U3314 ( .A(n1182), .B(n4385), .S0(n4330), .Y(n2474) );
  MXI2X1 U3315 ( .A(n1181), .B(n4386), .S0(n4330), .Y(n2476) );
  MXI2X1 U3316 ( .A(n1180), .B(n4383), .S0(n4330), .Y(n2478) );
  MXI2X1 U3317 ( .A(n1179), .B(n4384), .S0(n4330), .Y(n2480) );
  MXI2X1 U3318 ( .A(n1178), .B(n4381), .S0(n4330), .Y(n2482) );
  MXI2X1 U3319 ( .A(n1177), .B(n4382), .S0(n4330), .Y(n2484) );
  MXI2X1 U3320 ( .A(n1176), .B(n4379), .S0(n4330), .Y(n2486) );
  MXI2X1 U3321 ( .A(n1175), .B(n4380), .S0(n4330), .Y(n2488) );
  MXI2X1 U3322 ( .A(n1174), .B(n4377), .S0(n4330), .Y(n2490) );
  MXI2X1 U3323 ( .A(n1173), .B(n4378), .S0(n4330), .Y(n2492) );
  MXI2X1 U3324 ( .A(n1172), .B(n4375), .S0(n4329), .Y(n2494) );
  MXI2X1 U3325 ( .A(n1171), .B(n4376), .S0(n4330), .Y(n2496) );
  MXI2X1 U3326 ( .A(n1170), .B(n4373), .S0(n128), .Y(n2498) );
  MXI2X1 U3327 ( .A(n1169), .B(n4701), .S0(n128), .Y(n2500) );
  MXI2X1 U3328 ( .A(n1168), .B(n4670), .S0(n128), .Y(n2502) );
  MXI2X1 U3329 ( .A(n1167), .B(n4372), .S0(n128), .Y(n2504) );
  MXI2X1 U3330 ( .A(n1166), .B(n4369), .S0(n128), .Y(n2506) );
  MXI2X1 U3331 ( .A(n1165), .B(n4370), .S0(n128), .Y(n2508) );
  MXI2X1 U3332 ( .A(n1164), .B(n4952), .S0(n4331), .Y(n2510) );
  MXI2X1 U3333 ( .A(n1163), .B(n4966), .S0(n4331), .Y(n2512) );
  MXI2X1 U3334 ( .A(n1162), .B(n4934), .S0(n4331), .Y(n2514) );
  MXI2X1 U3335 ( .A(n1161), .B(n4943), .S0(n4331), .Y(n2516) );
  MXI2X1 U3336 ( .A(n1160), .B(n4913), .S0(n4331), .Y(n2518) );
  MXI2X1 U3337 ( .A(n1159), .B(n4922), .S0(n4331), .Y(n2520) );
  MXI2X1 U3338 ( .A(n1158), .B(n4895), .S0(n4331), .Y(n2522) );
  MXI2X1 U3339 ( .A(n1157), .B(n4904), .S0(n4331), .Y(n2524) );
  MXI2X1 U3340 ( .A(n1156), .B(n4874), .S0(n4331), .Y(n2526) );
  MXI2X1 U3341 ( .A(n1155), .B(n4883), .S0(n4331), .Y(n2528) );
  MXI2X1 U3342 ( .A(n1154), .B(n4856), .S0(n4331), .Y(n2530) );
  MXI2X1 U3343 ( .A(n1153), .B(n4865), .S0(n4331), .Y(n2532) );
  MXI2X1 U3344 ( .A(n1152), .B(n4834), .S0(n4332), .Y(n2534) );
  MXI2X1 U3345 ( .A(n1151), .B(n4843), .S0(n4332), .Y(n2536) );
  MXI2X1 U3346 ( .A(n1150), .B(n4816), .S0(n4332), .Y(n2538) );
  MXI2X1 U3347 ( .A(n1149), .B(n4825), .S0(n4332), .Y(n2540) );
  MXI2X1 U3348 ( .A(n1148), .B(n4790), .S0(n4332), .Y(n2542) );
  MXI2X1 U3349 ( .A(n1147), .B(n4799), .S0(n4332), .Y(n2544) );
  MXI2X1 U3350 ( .A(n1146), .B(n4772), .S0(n4332), .Y(n2546) );
  MXI2X1 U3351 ( .A(n1145), .B(n4781), .S0(n4332), .Y(n2548) );
  MXI2X1 U3352 ( .A(n1144), .B(n4750), .S0(n4332), .Y(n2550) );
  MXI2X1 U3353 ( .A(n1143), .B(n4759), .S0(n4332), .Y(n2552) );
  MXI2X1 U3354 ( .A(n1142), .B(n4732), .S0(n4332), .Y(n2554) );
  MXI2X1 U3355 ( .A(n1141), .B(n4741), .S0(n4332), .Y(n2556) );
  MXI2X1 U3356 ( .A(n1140), .B(n4710), .S0(n4331), .Y(n2558) );
  MXI2X1 U3357 ( .A(n1139), .B(n4719), .S0(n4332), .Y(n2560) );
  MXI2X1 U3358 ( .A(n1138), .B(n4692), .S0(n109), .Y(n2562) );
  MXI2X1 U3359 ( .A(n1137), .B(n4701), .S0(n109), .Y(n2564) );
  MXI2X1 U3360 ( .A(n1136), .B(n4670), .S0(n109), .Y(n2566) );
  MXI2X1 U3361 ( .A(n1135), .B(n4679), .S0(n109), .Y(n2568) );
  MXI2X1 U3362 ( .A(n1134), .B(n4652), .S0(n109), .Y(n2570) );
  MXI2X1 U3363 ( .A(n1133), .B(n4661), .S0(n109), .Y(n2572) );
  MXI2X1 U3364 ( .A(n1132), .B(n4952), .S0(n4333), .Y(n2574) );
  MXI2X1 U3365 ( .A(n1131), .B(n4966), .S0(n4333), .Y(n2576) );
  MXI2X1 U3366 ( .A(n1130), .B(n4934), .S0(n4333), .Y(n2578) );
  MXI2X1 U3367 ( .A(n1129), .B(n4943), .S0(n4333), .Y(n2580) );
  MXI2X1 U3368 ( .A(n1128), .B(n4913), .S0(n4333), .Y(n2582) );
  MXI2X1 U3369 ( .A(n1127), .B(n4922), .S0(n4333), .Y(n2584) );
  MXI2X1 U3370 ( .A(n1126), .B(n4895), .S0(n4333), .Y(n2586) );
  MXI2X1 U3371 ( .A(n1125), .B(n4904), .S0(n4333), .Y(n2588) );
  MXI2X1 U3372 ( .A(n1124), .B(n4874), .S0(n4333), .Y(n2590) );
  MXI2X1 U3373 ( .A(n1123), .B(n4883), .S0(n4333), .Y(n2592) );
  MXI2X1 U3374 ( .A(n1122), .B(n4856), .S0(n4333), .Y(n2594) );
  MXI2X1 U3375 ( .A(n1121), .B(n4865), .S0(n4333), .Y(n2596) );
  MXI2X1 U3376 ( .A(n1120), .B(n4834), .S0(n4334), .Y(n2598) );
  MXI2X1 U3377 ( .A(n1119), .B(n4843), .S0(n4334), .Y(n2600) );
  MXI2X1 U3378 ( .A(n1118), .B(n4816), .S0(n4334), .Y(n2602) );
  MXI2X1 U3379 ( .A(n1117), .B(n4825), .S0(n4334), .Y(n2604) );
  MXI2X1 U3380 ( .A(n1116), .B(n4790), .S0(n4334), .Y(n2606) );
  MXI2X1 U3381 ( .A(n1115), .B(n4799), .S0(n4334), .Y(n2608) );
  MXI2X1 U3382 ( .A(n1114), .B(n4772), .S0(n4334), .Y(n2610) );
  MXI2X1 U3383 ( .A(n1113), .B(n4781), .S0(n4334), .Y(n2612) );
  MXI2X1 U3384 ( .A(n1112), .B(n4750), .S0(n4334), .Y(n2614) );
  MXI2X1 U3385 ( .A(n1111), .B(n4759), .S0(n4334), .Y(n2616) );
  MXI2X1 U3386 ( .A(n1110), .B(n4732), .S0(n4334), .Y(n2618) );
  MXI2X1 U3387 ( .A(n1109), .B(n4741), .S0(n4334), .Y(n2620) );
  MXI2X1 U3388 ( .A(n1108), .B(n4710), .S0(n4333), .Y(n2622) );
  MXI2X1 U3389 ( .A(n1107), .B(n4719), .S0(n4334), .Y(n2624) );
  MXI2X1 U3390 ( .A(n1106), .B(n4692), .S0(n119), .Y(n2626) );
  MXI2X1 U3391 ( .A(n1105), .B(n4701), .S0(n119), .Y(n2628) );
  MXI2X1 U3392 ( .A(n1104), .B(n4670), .S0(n119), .Y(n2630) );
  MXI2X1 U3393 ( .A(n1103), .B(n4679), .S0(n119), .Y(n2632) );
  MXI2X1 U3394 ( .A(n1102), .B(n4652), .S0(n119), .Y(n2634) );
  MXI2X1 U3395 ( .A(n1101), .B(n4661), .S0(n119), .Y(n2636) );
  MXI2X1 U3396 ( .A(n1100), .B(n4952), .S0(n4335), .Y(n2638) );
  MXI2X1 U3397 ( .A(n1099), .B(n4966), .S0(n4335), .Y(n2640) );
  MXI2X1 U3398 ( .A(n1098), .B(n4934), .S0(n4335), .Y(n2642) );
  MXI2X1 U3399 ( .A(n1097), .B(n4943), .S0(n4335), .Y(n2644) );
  MXI2X1 U3400 ( .A(n1096), .B(n4913), .S0(n4335), .Y(n2646) );
  MXI2X1 U3401 ( .A(n1095), .B(n4922), .S0(n4335), .Y(n2648) );
  MXI2X1 U3402 ( .A(n1094), .B(n4895), .S0(n4335), .Y(n2650) );
  MXI2X1 U3403 ( .A(n1093), .B(n4904), .S0(n4335), .Y(n2652) );
  MXI2X1 U3404 ( .A(n1092), .B(n4874), .S0(n4335), .Y(n2654) );
  MXI2X1 U3405 ( .A(n1091), .B(n4883), .S0(n4335), .Y(n2656) );
  MXI2X1 U3406 ( .A(n1090), .B(n4856), .S0(n4335), .Y(n2658) );
  MXI2X1 U3407 ( .A(n1089), .B(n4865), .S0(n4335), .Y(n2660) );
  MXI2X1 U3408 ( .A(n1088), .B(n4834), .S0(n4336), .Y(n2662) );
  MXI2X1 U3409 ( .A(n1087), .B(n4843), .S0(n4336), .Y(n2664) );
  MXI2X1 U3410 ( .A(n1086), .B(n4816), .S0(n4336), .Y(n2666) );
  MXI2X1 U3411 ( .A(n1085), .B(n4825), .S0(n4336), .Y(n2668) );
  MXI2X1 U3412 ( .A(n1084), .B(n4790), .S0(n4336), .Y(n2670) );
  MXI2X1 U3413 ( .A(n1083), .B(n4799), .S0(n4336), .Y(n2672) );
  MXI2X1 U3414 ( .A(n1082), .B(n4772), .S0(n4336), .Y(n2674) );
  MXI2X1 U3415 ( .A(n1081), .B(n4781), .S0(n4336), .Y(n2676) );
  MXI2X1 U3416 ( .A(n1080), .B(n4750), .S0(n4336), .Y(n2678) );
  MXI2X1 U3417 ( .A(n1079), .B(n4759), .S0(n4336), .Y(n2680) );
  MXI2X1 U3418 ( .A(n1078), .B(n4732), .S0(n4336), .Y(n2682) );
  MXI2X1 U3419 ( .A(n1077), .B(n4741), .S0(n4336), .Y(n2684) );
  MXI2X1 U3420 ( .A(n1076), .B(n4710), .S0(n4335), .Y(n2686) );
  MXI2X1 U3421 ( .A(n1075), .B(n4719), .S0(n4336), .Y(n2688) );
  MXI2X1 U3422 ( .A(n1074), .B(n4692), .S0(n138), .Y(n2690) );
  MXI2X1 U3423 ( .A(n1073), .B(n4701), .S0(n138), .Y(n2692) );
  MXI2X1 U3424 ( .A(n1072), .B(n4670), .S0(n138), .Y(n2694) );
  MXI2X1 U3425 ( .A(n1071), .B(n4679), .S0(n138), .Y(n2696) );
  MXI2X1 U3426 ( .A(n1070), .B(n4652), .S0(n138), .Y(n2698) );
  MXI2X1 U3427 ( .A(n1069), .B(n4661), .S0(n138), .Y(n2700) );
  MXI2X1 U3428 ( .A(n1068), .B(n4952), .S0(n4337), .Y(n2702) );
  MXI2X1 U3429 ( .A(n1067), .B(n4966), .S0(n4337), .Y(n2704) );
  MXI2X1 U3430 ( .A(n1066), .B(n4934), .S0(n4337), .Y(n2706) );
  MXI2X1 U3431 ( .A(n1065), .B(n4943), .S0(n4337), .Y(n2708) );
  MXI2X1 U3432 ( .A(n1064), .B(n4913), .S0(n4337), .Y(n2710) );
  MXI2X1 U3433 ( .A(n1063), .B(n4922), .S0(n4337), .Y(n2712) );
  MXI2X1 U3434 ( .A(n1062), .B(n4895), .S0(n4337), .Y(n2714) );
  MXI2X1 U3435 ( .A(n1061), .B(n4904), .S0(n4337), .Y(n2716) );
  MXI2X1 U3436 ( .A(n1060), .B(n4874), .S0(n4337), .Y(n2718) );
  MXI2X1 U3437 ( .A(n1059), .B(n4883), .S0(n4337), .Y(n2720) );
  MXI2X1 U3438 ( .A(n1058), .B(n4856), .S0(n4337), .Y(n2722) );
  MXI2X1 U3439 ( .A(n1057), .B(n4865), .S0(n4337), .Y(n2724) );
  MXI2X1 U3440 ( .A(n1056), .B(n4834), .S0(n4338), .Y(n2726) );
  MXI2X1 U3441 ( .A(n1055), .B(n4843), .S0(n4338), .Y(n2728) );
  MXI2X1 U3442 ( .A(n1054), .B(n4816), .S0(n4338), .Y(n2730) );
  MXI2X1 U3443 ( .A(n1053), .B(n4825), .S0(n4338), .Y(n2732) );
  MXI2X1 U3444 ( .A(n1052), .B(n4790), .S0(n4338), .Y(n2734) );
  MXI2X1 U3445 ( .A(n1051), .B(n4799), .S0(n4338), .Y(n2736) );
  MXI2X1 U3446 ( .A(n1050), .B(n4772), .S0(n4338), .Y(n2738) );
  MXI2X1 U3447 ( .A(n1049), .B(n4781), .S0(n4338), .Y(n2740) );
  MXI2X1 U3448 ( .A(n1048), .B(n4750), .S0(n4338), .Y(n2742) );
  MXI2X1 U3449 ( .A(n1047), .B(n4759), .S0(n4338), .Y(n2744) );
  MXI2X1 U3450 ( .A(n1046), .B(n4732), .S0(n4338), .Y(n2746) );
  MXI2X1 U3451 ( .A(n1045), .B(n4741), .S0(n4338), .Y(n2748) );
  MXI2X1 U3452 ( .A(n1044), .B(n4710), .S0(n4337), .Y(n2750) );
  MXI2X1 U3453 ( .A(n1043), .B(n4719), .S0(n4338), .Y(n2752) );
  MXI2X1 U3454 ( .A(n1042), .B(n4692), .S0(n129), .Y(n2754) );
  MXI2X1 U3455 ( .A(n1041), .B(n4701), .S0(n129), .Y(n2756) );
  MXI2X1 U3456 ( .A(n1040), .B(n4670), .S0(n129), .Y(n2758) );
  MXI2X1 U3457 ( .A(n1039), .B(n4679), .S0(n129), .Y(n2760) );
  MXI2X1 U3458 ( .A(n1038), .B(n4652), .S0(n129), .Y(n2762) );
  MXI2X1 U3459 ( .A(n1037), .B(n4661), .S0(n129), .Y(n2764) );
  MXI2X1 U3460 ( .A(n1036), .B(n4952), .S0(n4339), .Y(n2766) );
  MXI2X1 U3461 ( .A(n1035), .B(n4966), .S0(n4339), .Y(n2768) );
  MXI2X1 U3462 ( .A(n1034), .B(n4934), .S0(n4339), .Y(n2770) );
  MXI2X1 U3463 ( .A(n1033), .B(n4943), .S0(n4339), .Y(n2772) );
  MXI2X1 U3464 ( .A(n1032), .B(n4913), .S0(n4339), .Y(n2774) );
  MXI2X1 U3465 ( .A(n1031), .B(n4922), .S0(n4339), .Y(n2776) );
  MXI2X1 U3466 ( .A(n1030), .B(n4895), .S0(n4339), .Y(n2778) );
  MXI2X1 U3467 ( .A(n1029), .B(n4904), .S0(n4339), .Y(n2780) );
  MXI2X1 U3468 ( .A(n1028), .B(n4874), .S0(n4339), .Y(n2782) );
  MXI2X1 U3469 ( .A(n1027), .B(n4883), .S0(n4339), .Y(n2784) );
  MXI2X1 U3470 ( .A(n1026), .B(n4856), .S0(n4339), .Y(n2786) );
  MXI2X1 U3471 ( .A(n1025), .B(n4865), .S0(n4339), .Y(n2788) );
  MXI2X1 U3472 ( .A(n1024), .B(n4834), .S0(n4340), .Y(n2790) );
  MXI2X1 U3473 ( .A(n1023), .B(n4843), .S0(n4340), .Y(n2792) );
  MXI2X1 U3474 ( .A(n1022), .B(n4816), .S0(n4340), .Y(n2794) );
  MXI2X1 U3475 ( .A(n1021), .B(n4825), .S0(n4340), .Y(n2796) );
  MXI2X1 U3476 ( .A(n1020), .B(n4790), .S0(n4340), .Y(n2798) );
  MXI2X1 U3477 ( .A(n1019), .B(n4799), .S0(n4340), .Y(n2800) );
  MXI2X1 U3478 ( .A(n1018), .B(n4772), .S0(n4340), .Y(n2802) );
  MXI2X1 U3479 ( .A(n1017), .B(n4781), .S0(n4340), .Y(n2804) );
  MXI2X1 U3480 ( .A(n1016), .B(n4750), .S0(n4340), .Y(n2806) );
  MXI2X1 U3481 ( .A(n1015), .B(n4759), .S0(n4340), .Y(n2808) );
  MXI2X1 U3482 ( .A(n1014), .B(n4732), .S0(n4340), .Y(n2810) );
  MXI2X1 U3483 ( .A(n1013), .B(n4741), .S0(n4340), .Y(n2812) );
  MXI2X1 U3484 ( .A(n1012), .B(n4710), .S0(n4339), .Y(n2814) );
  MXI2X1 U3485 ( .A(n1011), .B(n4719), .S0(n4340), .Y(n2816) );
  MXI2X1 U3486 ( .A(n1010), .B(n4692), .S0(n110), .Y(n2818) );
  MXI2X1 U3487 ( .A(n1009), .B(n4701), .S0(n110), .Y(n2820) );
  MXI2X1 U3488 ( .A(n1008), .B(n4670), .S0(n110), .Y(n2822) );
  MXI2X1 U3489 ( .A(n1007), .B(n4679), .S0(n110), .Y(n2824) );
  MXI2X1 U3490 ( .A(n1006), .B(n4652), .S0(n110), .Y(n2826) );
  MXI2X1 U3491 ( .A(n1005), .B(n4661), .S0(n110), .Y(n2828) );
  MXI2X1 U3492 ( .A(n1004), .B(n4952), .S0(n4341), .Y(n2830) );
  MXI2X1 U3493 ( .A(n1003), .B(n4966), .S0(n4341), .Y(n2832) );
  MXI2X1 U3494 ( .A(n1002), .B(n4934), .S0(n4341), .Y(n2834) );
  MXI2X1 U3495 ( .A(n1001), .B(n4943), .S0(n4341), .Y(n2836) );
  MXI2X1 U3496 ( .A(n1000), .B(n4913), .S0(n4341), .Y(n2838) );
  MXI2X1 U3497 ( .A(n999), .B(n4922), .S0(n4341), .Y(n2840) );
  MXI2X1 U3498 ( .A(n998), .B(n4895), .S0(n4341), .Y(n2842) );
  MXI2X1 U3499 ( .A(n997), .B(n4904), .S0(n4341), .Y(n2844) );
  MXI2X1 U3500 ( .A(n996), .B(n4874), .S0(n4341), .Y(n2846) );
  MXI2X1 U3501 ( .A(n995), .B(n4883), .S0(n4341), .Y(n2848) );
  MXI2X1 U3502 ( .A(n994), .B(n4856), .S0(n4341), .Y(n2850) );
  MXI2X1 U3503 ( .A(n993), .B(n4865), .S0(n4341), .Y(n2852) );
  MXI2X1 U3504 ( .A(n992), .B(n4834), .S0(n4342), .Y(n2854) );
  MXI2X1 U3505 ( .A(n991), .B(n4843), .S0(n4342), .Y(n2856) );
  MXI2X1 U3506 ( .A(n990), .B(n4816), .S0(n4342), .Y(n2858) );
  MXI2X1 U3507 ( .A(n989), .B(n4825), .S0(n4342), .Y(n2860) );
  MXI2X1 U3508 ( .A(n988), .B(n4790), .S0(n4342), .Y(n2862) );
  MXI2X1 U3509 ( .A(n987), .B(n4799), .S0(n4342), .Y(n2864) );
  MXI2X1 U3510 ( .A(n986), .B(n4772), .S0(n4342), .Y(n2866) );
  MXI2X1 U3511 ( .A(n985), .B(n4781), .S0(n4342), .Y(n2868) );
  MXI2X1 U3512 ( .A(n984), .B(n4750), .S0(n4342), .Y(n2870) );
  MXI2X1 U3513 ( .A(n983), .B(n4759), .S0(n4342), .Y(n2872) );
  MXI2X1 U3514 ( .A(n982), .B(n4732), .S0(n4342), .Y(n2874) );
  MXI2X1 U3515 ( .A(n981), .B(n4741), .S0(n4342), .Y(n2876) );
  MXI2X1 U3516 ( .A(n980), .B(n4710), .S0(n4341), .Y(n2878) );
  MXI2X1 U3517 ( .A(n979), .B(n4719), .S0(n4342), .Y(n2880) );
  MXI2X1 U3518 ( .A(n978), .B(n4692), .S0(n120), .Y(n2882) );
  MXI2X1 U3519 ( .A(n977), .B(n4701), .S0(n120), .Y(n2884) );
  MXI2X1 U3520 ( .A(n976), .B(n4670), .S0(n120), .Y(n2886) );
  MXI2X1 U3521 ( .A(n975), .B(n4679), .S0(n120), .Y(n2888) );
  MXI2X1 U3522 ( .A(n974), .B(n4652), .S0(n120), .Y(n2890) );
  MXI2X1 U3523 ( .A(n973), .B(n4661), .S0(n120), .Y(n2892) );
  MXI2X1 U3524 ( .A(n972), .B(n4952), .S0(n4343), .Y(n2894) );
  MXI2X1 U3525 ( .A(n971), .B(n4966), .S0(n4343), .Y(n2896) );
  MXI2X1 U3526 ( .A(n970), .B(n4934), .S0(n4343), .Y(n2898) );
  MXI2X1 U3527 ( .A(n969), .B(n4943), .S0(n4343), .Y(n2900) );
  MXI2X1 U3528 ( .A(n968), .B(n4913), .S0(n4343), .Y(n2902) );
  MXI2X1 U3529 ( .A(n967), .B(n4922), .S0(n4343), .Y(n2904) );
  MXI2X1 U3530 ( .A(n966), .B(n4895), .S0(n4343), .Y(n2906) );
  MXI2X1 U3531 ( .A(n965), .B(n4904), .S0(n4343), .Y(n2908) );
  MXI2X1 U3532 ( .A(n964), .B(n4874), .S0(n4343), .Y(n2910) );
  MXI2X1 U3533 ( .A(n963), .B(n4883), .S0(n4343), .Y(n2912) );
  MXI2X1 U3534 ( .A(n962), .B(n4856), .S0(n4343), .Y(n2914) );
  MXI2X1 U3535 ( .A(n961), .B(n4865), .S0(n4343), .Y(n2916) );
  MXI2X1 U3536 ( .A(n960), .B(n4834), .S0(n4344), .Y(n2918) );
  MXI2X1 U3537 ( .A(n959), .B(n4843), .S0(n4344), .Y(n2920) );
  MXI2X1 U3538 ( .A(n958), .B(n4816), .S0(n4344), .Y(n2922) );
  MXI2X1 U3539 ( .A(n957), .B(n4825), .S0(n4344), .Y(n2924) );
  MXI2X1 U3540 ( .A(n956), .B(n4790), .S0(n4344), .Y(n2926) );
  MXI2X1 U3541 ( .A(n955), .B(n4799), .S0(n4344), .Y(n2928) );
  MXI2X1 U3542 ( .A(n954), .B(n4772), .S0(n4344), .Y(n2930) );
  MXI2X1 U3543 ( .A(n953), .B(n4781), .S0(n4344), .Y(n2932) );
  MXI2X1 U3544 ( .A(n952), .B(n4750), .S0(n4344), .Y(n2934) );
  MXI2X1 U3545 ( .A(n951), .B(n4759), .S0(n4344), .Y(n2936) );
  MXI2X1 U3546 ( .A(n950), .B(n4732), .S0(n4344), .Y(n2938) );
  MXI2X1 U3547 ( .A(n949), .B(n4741), .S0(n4344), .Y(n2940) );
  MXI2X1 U3548 ( .A(n948), .B(n4710), .S0(n4343), .Y(n2942) );
  MXI2X1 U3549 ( .A(n947), .B(n4719), .S0(n4344), .Y(n2944) );
  MXI2X1 U3550 ( .A(n946), .B(n4692), .S0(n139), .Y(n2946) );
  MXI2X1 U3551 ( .A(n945), .B(n4701), .S0(n139), .Y(n2948) );
  MXI2X1 U3552 ( .A(n944), .B(n4670), .S0(n139), .Y(n2950) );
  MXI2X1 U3553 ( .A(n943), .B(n4679), .S0(n139), .Y(n2952) );
  MXI2X1 U3554 ( .A(n942), .B(n4652), .S0(n139), .Y(n2954) );
  MXI2X1 U3555 ( .A(n941), .B(n4661), .S0(n139), .Y(n2956) );
  MXI2X1 U3556 ( .A(n940), .B(n4952), .S0(n4345), .Y(n2958) );
  MXI2X1 U3557 ( .A(n939), .B(n4966), .S0(n4345), .Y(n2960) );
  MXI2X1 U3558 ( .A(n938), .B(n4934), .S0(n4345), .Y(n2962) );
  MXI2X1 U3559 ( .A(n937), .B(n4943), .S0(n4345), .Y(n2964) );
  MXI2X1 U3560 ( .A(n936), .B(n4913), .S0(n4345), .Y(n2966) );
  MXI2X1 U3561 ( .A(n935), .B(n4922), .S0(n4345), .Y(n2968) );
  MXI2X1 U3562 ( .A(n934), .B(n4895), .S0(n4345), .Y(n2970) );
  MXI2X1 U3563 ( .A(n933), .B(n4904), .S0(n4345), .Y(n2972) );
  MXI2X1 U3564 ( .A(n932), .B(n4874), .S0(n4345), .Y(n2974) );
  MXI2X1 U3565 ( .A(n931), .B(n4883), .S0(n4345), .Y(n2976) );
  MXI2X1 U3566 ( .A(n930), .B(n4856), .S0(n4345), .Y(n2978) );
  MXI2X1 U3567 ( .A(n929), .B(n4865), .S0(n4345), .Y(n2980) );
  MXI2X1 U3568 ( .A(n928), .B(n4834), .S0(n4346), .Y(n2982) );
  MXI2X1 U3569 ( .A(n927), .B(n4843), .S0(n4346), .Y(n2984) );
  MXI2X1 U3570 ( .A(n926), .B(n4816), .S0(n4346), .Y(n2986) );
  MXI2X1 U3571 ( .A(n925), .B(n4825), .S0(n4346), .Y(n2988) );
  MXI2X1 U3572 ( .A(n924), .B(n4790), .S0(n4346), .Y(n2990) );
  MXI2X1 U3573 ( .A(n923), .B(n4799), .S0(n4346), .Y(n2992) );
  MXI2X1 U3574 ( .A(n922), .B(n4772), .S0(n4346), .Y(n2994) );
  MXI2X1 U3575 ( .A(n921), .B(n4781), .S0(n4346), .Y(n2996) );
  MXI2X1 U3576 ( .A(n920), .B(n4750), .S0(n4346), .Y(n2998) );
  MXI2X1 U3577 ( .A(n919), .B(n4759), .S0(n4346), .Y(n3000) );
  MXI2X1 U3578 ( .A(n918), .B(n4732), .S0(n4346), .Y(n3002) );
  MXI2X1 U3579 ( .A(n917), .B(n4741), .S0(n4346), .Y(n3004) );
  MXI2X1 U3580 ( .A(n916), .B(n4710), .S0(n4345), .Y(n3006) );
  MXI2X1 U3581 ( .A(n915), .B(n4719), .S0(n4346), .Y(n3008) );
  MXI2X1 U3582 ( .A(n914), .B(n4692), .S0(n130), .Y(n3010) );
  MXI2X1 U3583 ( .A(n913), .B(n4701), .S0(n130), .Y(n3012) );
  MXI2X1 U3584 ( .A(n912), .B(n4670), .S0(n130), .Y(n3014) );
  MXI2X1 U3585 ( .A(n911), .B(n4679), .S0(n130), .Y(n3016) );
  MXI2X1 U3586 ( .A(n910), .B(n4652), .S0(n130), .Y(n3018) );
  MXI2X1 U3587 ( .A(n909), .B(n4661), .S0(n130), .Y(n3020) );
  MXI2X1 U3588 ( .A(n908), .B(n4952), .S0(n4347), .Y(n3022) );
  MXI2X1 U3589 ( .A(n907), .B(n4966), .S0(n4347), .Y(n3024) );
  MXI2X1 U3590 ( .A(n906), .B(n4934), .S0(n4347), .Y(n3026) );
  MXI2X1 U3591 ( .A(n905), .B(n4943), .S0(n4347), .Y(n3028) );
  MXI2X1 U3592 ( .A(n904), .B(n4913), .S0(n4347), .Y(n3030) );
  MXI2X1 U3593 ( .A(n903), .B(n4922), .S0(n4347), .Y(n3032) );
  MXI2X1 U3594 ( .A(n902), .B(n4895), .S0(n4347), .Y(n3034) );
  MXI2X1 U3595 ( .A(n901), .B(n4904), .S0(n4347), .Y(n3036) );
  MXI2X1 U3596 ( .A(n900), .B(n4874), .S0(n4347), .Y(n3038) );
  MXI2X1 U3597 ( .A(n899), .B(n4883), .S0(n4347), .Y(n3040) );
  MXI2X1 U3598 ( .A(n898), .B(n4856), .S0(n4347), .Y(n3042) );
  MXI2X1 U3599 ( .A(n897), .B(n4865), .S0(n4347), .Y(n3044) );
  MXI2X1 U3600 ( .A(n896), .B(n4834), .S0(n4348), .Y(n3046) );
  MXI2X1 U3601 ( .A(n895), .B(n4843), .S0(n4348), .Y(n3048) );
  MXI2X1 U3602 ( .A(n894), .B(n4816), .S0(n4348), .Y(n3050) );
  MXI2X1 U3603 ( .A(n893), .B(n4825), .S0(n4348), .Y(n3052) );
  MXI2X1 U3604 ( .A(n892), .B(n4790), .S0(n4348), .Y(n3054) );
  MXI2X1 U3605 ( .A(n891), .B(n4799), .S0(n4348), .Y(n3056) );
  MXI2X1 U3606 ( .A(n890), .B(n4772), .S0(n4348), .Y(n3058) );
  MXI2X1 U3607 ( .A(n889), .B(n4781), .S0(n4348), .Y(n3060) );
  MXI2X1 U3608 ( .A(n888), .B(n4750), .S0(n4348), .Y(n3062) );
  MXI2X1 U3609 ( .A(n887), .B(n4759), .S0(n4348), .Y(n3064) );
  MXI2X1 U3610 ( .A(n886), .B(n4732), .S0(n4348), .Y(n3066) );
  MXI2X1 U3611 ( .A(n885), .B(n4741), .S0(n4348), .Y(n3068) );
  MXI2X1 U3612 ( .A(n884), .B(n4710), .S0(n4347), .Y(n3070) );
  MXI2X1 U3613 ( .A(n883), .B(n4719), .S0(n4348), .Y(n3072) );
  MXI2X1 U3614 ( .A(n882), .B(n4692), .S0(n111), .Y(n3074) );
  MXI2X1 U3615 ( .A(n881), .B(n4701), .S0(n111), .Y(n3076) );
  MXI2X1 U3616 ( .A(n880), .B(n4670), .S0(n111), .Y(n3078) );
  MXI2X1 U3617 ( .A(n879), .B(n4679), .S0(n111), .Y(n3080) );
  MXI2X1 U3618 ( .A(n878), .B(n4652), .S0(n111), .Y(n3082) );
  MXI2X1 U3619 ( .A(n877), .B(n4661), .S0(n111), .Y(n3084) );
  MXI2X1 U3620 ( .A(n876), .B(n4952), .S0(n4349), .Y(n3086) );
  MXI2X1 U3621 ( .A(n875), .B(n4966), .S0(n4349), .Y(n3088) );
  MXI2X1 U3622 ( .A(n874), .B(n4934), .S0(n4349), .Y(n3090) );
  MXI2X1 U3623 ( .A(n873), .B(n4943), .S0(n4349), .Y(n3092) );
  MXI2X1 U3624 ( .A(n872), .B(n4913), .S0(n4349), .Y(n3094) );
  MXI2X1 U3625 ( .A(n871), .B(n4922), .S0(n4349), .Y(n3096) );
  MXI2X1 U3626 ( .A(n870), .B(n4895), .S0(n4349), .Y(n3098) );
  MXI2X1 U3627 ( .A(n869), .B(n4904), .S0(n4349), .Y(n3100) );
  MXI2X1 U3628 ( .A(n868), .B(n4874), .S0(n4349), .Y(n3102) );
  MXI2X1 U3629 ( .A(n867), .B(n4883), .S0(n4349), .Y(n3104) );
  MXI2X1 U3630 ( .A(n866), .B(n4856), .S0(n4349), .Y(n3106) );
  MXI2X1 U3631 ( .A(n865), .B(n4865), .S0(n4349), .Y(n3108) );
  MXI2X1 U3632 ( .A(n864), .B(n4834), .S0(n4350), .Y(n3110) );
  MXI2X1 U3633 ( .A(n863), .B(n4843), .S0(n4350), .Y(n3112) );
  MXI2X1 U3634 ( .A(n862), .B(n4816), .S0(n4350), .Y(n3114) );
  MXI2X1 U3635 ( .A(n861), .B(n4825), .S0(n4350), .Y(n3116) );
  MXI2X1 U3636 ( .A(n860), .B(n4790), .S0(n4350), .Y(n3118) );
  MXI2X1 U3637 ( .A(n859), .B(n4799), .S0(n4350), .Y(n3120) );
  MXI2X1 U3638 ( .A(n858), .B(n4772), .S0(n4350), .Y(n3122) );
  MXI2X1 U3639 ( .A(n857), .B(n4781), .S0(n4350), .Y(n3124) );
  MXI2X1 U3640 ( .A(n856), .B(n4750), .S0(n4350), .Y(n3126) );
  MXI2X1 U3641 ( .A(n855), .B(n4759), .S0(n4350), .Y(n3128) );
  MXI2X1 U3642 ( .A(n854), .B(n4732), .S0(n4350), .Y(n3130) );
  MXI2X1 U3643 ( .A(n853), .B(n4741), .S0(n4350), .Y(n3132) );
  MXI2X1 U3644 ( .A(n852), .B(n4710), .S0(n4349), .Y(n3134) );
  MXI2X1 U3645 ( .A(n851), .B(n4719), .S0(n4350), .Y(n3136) );
  MXI2X1 U3646 ( .A(n850), .B(n4692), .S0(n121), .Y(n3138) );
  MXI2X1 U3647 ( .A(n849), .B(n4701), .S0(n121), .Y(n3140) );
  MXI2X1 U3648 ( .A(n848), .B(n4670), .S0(n121), .Y(n3142) );
  MXI2X1 U3649 ( .A(n847), .B(n4679), .S0(n121), .Y(n3144) );
  MXI2X1 U3650 ( .A(n846), .B(n4652), .S0(n121), .Y(n3146) );
  MXI2X1 U3651 ( .A(n845), .B(n4661), .S0(n121), .Y(n3148) );
  MXI2X1 U3652 ( .A(n844), .B(n4952), .S0(n4351), .Y(n3150) );
  MXI2X1 U3653 ( .A(n843), .B(n4966), .S0(n4351), .Y(n3152) );
  MXI2X1 U3654 ( .A(n842), .B(n4934), .S0(n4351), .Y(n3154) );
  MXI2X1 U3655 ( .A(n841), .B(n4943), .S0(n4351), .Y(n3156) );
  MXI2X1 U3656 ( .A(n840), .B(n4913), .S0(n4351), .Y(n3158) );
  MXI2X1 U3657 ( .A(n839), .B(n4922), .S0(n4351), .Y(n3160) );
  MXI2X1 U3658 ( .A(n838), .B(n4895), .S0(n4351), .Y(n3162) );
  MXI2X1 U3659 ( .A(n837), .B(n4904), .S0(n4351), .Y(n3164) );
  MXI2X1 U3660 ( .A(n836), .B(n4874), .S0(n4351), .Y(n3166) );
  MXI2X1 U3661 ( .A(n835), .B(n4883), .S0(n4351), .Y(n3168) );
  MXI2X1 U3662 ( .A(n834), .B(n4856), .S0(n4351), .Y(n3170) );
  MXI2X1 U3663 ( .A(n833), .B(n4865), .S0(n4351), .Y(n3172) );
  MXI2X1 U3664 ( .A(n832), .B(n4834), .S0(n4352), .Y(n3174) );
  MXI2X1 U3665 ( .A(n831), .B(n4843), .S0(n4352), .Y(n3176) );
  MXI2X1 U3666 ( .A(n830), .B(n4816), .S0(n4352), .Y(n3178) );
  MXI2X1 U3667 ( .A(n829), .B(n4825), .S0(n4352), .Y(n3180) );
  MXI2X1 U3668 ( .A(n828), .B(n4790), .S0(n4352), .Y(n3182) );
  MXI2X1 U3669 ( .A(n827), .B(n4799), .S0(n4352), .Y(n3184) );
  MXI2X1 U3670 ( .A(n826), .B(n4772), .S0(n4352), .Y(n3186) );
  MXI2X1 U3671 ( .A(n825), .B(n4781), .S0(n4352), .Y(n3188) );
  MXI2X1 U3672 ( .A(n824), .B(n4750), .S0(n4352), .Y(n3190) );
  MXI2X1 U3673 ( .A(n823), .B(n4759), .S0(n4352), .Y(n3192) );
  MXI2X1 U3674 ( .A(n822), .B(n4732), .S0(n4352), .Y(n3194) );
  MXI2X1 U3675 ( .A(n821), .B(n4741), .S0(n4352), .Y(n3196) );
  MXI2X1 U3676 ( .A(n820), .B(n4710), .S0(n4351), .Y(n3198) );
  MXI2X1 U3677 ( .A(n819), .B(n4719), .S0(n4352), .Y(n3200) );
  MXI2X1 U3678 ( .A(n818), .B(n4692), .S0(n140), .Y(n3202) );
  MXI2X1 U3679 ( .A(n817), .B(n4701), .S0(n140), .Y(n3204) );
  MXI2X1 U3680 ( .A(n816), .B(n4670), .S0(n140), .Y(n3206) );
  MXI2X1 U3681 ( .A(n815), .B(n4679), .S0(n140), .Y(n3208) );
  MXI2X1 U3682 ( .A(n814), .B(n4652), .S0(n140), .Y(n3210) );
  MXI2X1 U3683 ( .A(n813), .B(n4661), .S0(n140), .Y(n3212) );
  MXI2X1 U3684 ( .A(n812), .B(n4399), .S0(n4353), .Y(n3214) );
  MXI2X1 U3685 ( .A(n811), .B(n4966), .S0(n4353), .Y(n3216) );
  MXI2X1 U3686 ( .A(n810), .B(n4934), .S0(n4353), .Y(n3218) );
  MXI2X1 U3687 ( .A(n809), .B(n4943), .S0(n4353), .Y(n3220) );
  MXI2X1 U3688 ( .A(n808), .B(n4913), .S0(n4353), .Y(n3222) );
  MXI2X1 U3689 ( .A(n807), .B(n4922), .S0(n4353), .Y(n3224) );
  MXI2X1 U3690 ( .A(n806), .B(n4895), .S0(n4353), .Y(n3226) );
  MXI2X1 U3691 ( .A(n805), .B(n4904), .S0(n4353), .Y(n3228) );
  MXI2X1 U3692 ( .A(n804), .B(n4874), .S0(n4353), .Y(n3230) );
  MXI2X1 U3693 ( .A(n803), .B(n4883), .S0(n4353), .Y(n3232) );
  MXI2X1 U3694 ( .A(n802), .B(n4856), .S0(n4353), .Y(n3234) );
  MXI2X1 U3695 ( .A(n801), .B(n4390), .S0(n4353), .Y(n3236) );
  MXI2X1 U3696 ( .A(n800), .B(n4834), .S0(n4354), .Y(n3238) );
  MXI2X1 U3697 ( .A(n799), .B(n4388), .S0(n4354), .Y(n3240) );
  MXI2X1 U3698 ( .A(n798), .B(n4816), .S0(n4354), .Y(n3242) );
  MXI2X1 U3699 ( .A(n797), .B(n4825), .S0(n4354), .Y(n3244) );
  MXI2X1 U3700 ( .A(n796), .B(n4383), .S0(n4354), .Y(n3246) );
  MXI2X1 U3701 ( .A(n795), .B(n4384), .S0(n4354), .Y(n3248) );
  MXI2X1 U3702 ( .A(n794), .B(n4381), .S0(n4354), .Y(n3250) );
  MXI2X1 U3703 ( .A(n793), .B(n4382), .S0(n4354), .Y(n3252) );
  MXI2X1 U3704 ( .A(n792), .B(n4379), .S0(n4354), .Y(n3254) );
  MXI2X1 U3705 ( .A(n791), .B(n4380), .S0(n4354), .Y(n3256) );
  MXI2X1 U3706 ( .A(n790), .B(n4377), .S0(n4354), .Y(n3258) );
  MXI2X1 U3707 ( .A(n789), .B(n4378), .S0(n4354), .Y(n3260) );
  MXI2X1 U3708 ( .A(n788), .B(n4710), .S0(n131), .Y(n3262) );
  MXI2X1 U3709 ( .A(n787), .B(n4719), .S0(n131), .Y(n3264) );
  MXI2X1 U3710 ( .A(n786), .B(n4692), .S0(n131), .Y(n3266) );
  MXI2X1 U3711 ( .A(n785), .B(n4374), .S0(n4353), .Y(n3268) );
  MXI2X1 U3712 ( .A(n784), .B(n4371), .S0(n4354), .Y(n3270) );
  MXI2X1 U3713 ( .A(n783), .B(n4372), .S0(n131), .Y(n3272) );
  MXI2X1 U3714 ( .A(n782), .B(n4369), .S0(n131), .Y(n3274) );
  MXI2X1 U3715 ( .A(n781), .B(n4370), .S0(n131), .Y(n3276) );
  MXI2X1 U3716 ( .A(n780), .B(n4952), .S0(n4355), .Y(n3278) );
  MXI2X1 U3717 ( .A(n779), .B(n4966), .S0(n4355), .Y(n3280) );
  MXI2X1 U3718 ( .A(n778), .B(n4934), .S0(n4355), .Y(n3282) );
  MXI2X1 U3719 ( .A(n777), .B(n4943), .S0(n4355), .Y(n3284) );
  MXI2X1 U3720 ( .A(n776), .B(n4913), .S0(n4355), .Y(n3286) );
  MXI2X1 U3721 ( .A(n775), .B(n4922), .S0(n4355), .Y(n3288) );
  MXI2X1 U3722 ( .A(n774), .B(n4895), .S0(n4355), .Y(n3290) );
  MXI2X1 U3723 ( .A(n773), .B(n4904), .S0(n4355), .Y(n3292) );
  MXI2X1 U3724 ( .A(n772), .B(n4874), .S0(n4355), .Y(n3294) );
  MXI2X1 U3725 ( .A(n771), .B(n4883), .S0(n4355), .Y(n3296) );
  MXI2X1 U3726 ( .A(n770), .B(n4856), .S0(n4355), .Y(n3298) );
  MXI2X1 U3727 ( .A(n769), .B(n4865), .S0(n4355), .Y(n3300) );
  MXI2X1 U3728 ( .A(n768), .B(n4834), .S0(n4356), .Y(n3302) );
  MXI2X1 U3729 ( .A(n767), .B(n4843), .S0(n4356), .Y(n3304) );
  MXI2X1 U3730 ( .A(n766), .B(n4816), .S0(n4356), .Y(n3306) );
  MXI2X1 U3731 ( .A(n765), .B(n4825), .S0(n4356), .Y(n3308) );
  MXI2X1 U3732 ( .A(n764), .B(n4790), .S0(n4356), .Y(n3310) );
  MXI2X1 U3733 ( .A(n763), .B(n4799), .S0(n4356), .Y(n3312) );
  MXI2X1 U3734 ( .A(n762), .B(n4772), .S0(n4356), .Y(n3314) );
  MXI2X1 U3735 ( .A(n761), .B(n4781), .S0(n4356), .Y(n3316) );
  MXI2X1 U3736 ( .A(n760), .B(n4750), .S0(n4356), .Y(n3318) );
  MXI2X1 U3737 ( .A(n759), .B(n4759), .S0(n4356), .Y(n3320) );
  MXI2X1 U3738 ( .A(n758), .B(n4732), .S0(n4356), .Y(n3322) );
  MXI2X1 U3739 ( .A(n757), .B(n4741), .S0(n4356), .Y(n3324) );
  MXI2X1 U3740 ( .A(n756), .B(n4710), .S0(n112), .Y(n3326) );
  MXI2X1 U3741 ( .A(n755), .B(n4719), .S0(n112), .Y(n3328) );
  MXI2X1 U3742 ( .A(n754), .B(n4692), .S0(n112), .Y(n3330) );
  MXI2X1 U3743 ( .A(n753), .B(n4374), .S0(n4355), .Y(n3332) );
  MXI2X1 U3744 ( .A(n752), .B(n4371), .S0(n4356), .Y(n3334) );
  MXI2X1 U3745 ( .A(n751), .B(n4679), .S0(n112), .Y(n3336) );
  MXI2X1 U3746 ( .A(n750), .B(n4652), .S0(n112), .Y(n3338) );
  MXI2X1 U3747 ( .A(n749), .B(n4661), .S0(n112), .Y(n3340) );
  MXI2X1 U3748 ( .A(n748), .B(n4952), .S0(n4357), .Y(n3342) );
  MXI2X1 U3749 ( .A(n747), .B(n4966), .S0(n4357), .Y(n3344) );
  MXI2X1 U3750 ( .A(n746), .B(n4934), .S0(n4357), .Y(n3346) );
  MXI2X1 U3751 ( .A(n745), .B(n4943), .S0(n4357), .Y(n3348) );
  MXI2X1 U3752 ( .A(n744), .B(n4913), .S0(n4357), .Y(n3350) );
  MXI2X1 U3753 ( .A(n743), .B(n4922), .S0(n4357), .Y(n3352) );
  MXI2X1 U3754 ( .A(n742), .B(n4895), .S0(n4357), .Y(n3354) );
  MXI2X1 U3755 ( .A(n741), .B(n4904), .S0(n4357), .Y(n3356) );
  MXI2X1 U3756 ( .A(n740), .B(n4874), .S0(n4357), .Y(n3358) );
  MXI2X1 U3757 ( .A(n739), .B(n4883), .S0(n4357), .Y(n3360) );
  MXI2X1 U3758 ( .A(n738), .B(n4856), .S0(n4357), .Y(n3362) );
  MXI2X1 U3759 ( .A(n737), .B(n4865), .S0(n4357), .Y(n3364) );
  MXI2X1 U3760 ( .A(n736), .B(n4834), .S0(n4358), .Y(n3366) );
  MXI2X1 U3761 ( .A(n735), .B(n4843), .S0(n4358), .Y(n3368) );
  MXI2X1 U3762 ( .A(n734), .B(n4816), .S0(n4358), .Y(n3370) );
  MXI2X1 U3763 ( .A(n733), .B(n4825), .S0(n4358), .Y(n3372) );
  MXI2X1 U3764 ( .A(n732), .B(n4790), .S0(n4358), .Y(n3374) );
  MXI2X1 U3765 ( .A(n731), .B(n4799), .S0(n4358), .Y(n3376) );
  MXI2X1 U3766 ( .A(n730), .B(n4772), .S0(n4358), .Y(n3378) );
  MXI2X1 U3767 ( .A(n729), .B(n4781), .S0(n4358), .Y(n3380) );
  MXI2X1 U3768 ( .A(n728), .B(n4750), .S0(n4358), .Y(n3382) );
  MXI2X1 U3769 ( .A(n727), .B(n4759), .S0(n4358), .Y(n3384) );
  MXI2X1 U3770 ( .A(n726), .B(n4732), .S0(n4358), .Y(n3386) );
  MXI2X1 U3771 ( .A(n725), .B(n4741), .S0(n4358), .Y(n3388) );
  MXI2X1 U3772 ( .A(n724), .B(n4710), .S0(n4357), .Y(n3390) );
  MXI2X1 U3773 ( .A(n723), .B(n4719), .S0(n4358), .Y(n3392) );
  MXI2X1 U3774 ( .A(n722), .B(n4692), .S0(n122), .Y(n3394) );
  MXI2X1 U3775 ( .A(n721), .B(n4701), .S0(n122), .Y(n3396) );
  MXI2X1 U3776 ( .A(n720), .B(n4670), .S0(n122), .Y(n3398) );
  MXI2X1 U3777 ( .A(n719), .B(n4679), .S0(n122), .Y(n3400) );
  MXI2X1 U3778 ( .A(n718), .B(n4652), .S0(n122), .Y(n3402) );
  MXI2X1 U3779 ( .A(n717), .B(n4661), .S0(n122), .Y(n3404) );
  MXI2X1 U3780 ( .A(n716), .B(n4952), .S0(n4359), .Y(n3406) );
  MXI2X1 U3781 ( .A(n715), .B(n4966), .S0(n4359), .Y(n3408) );
  MXI2X1 U3782 ( .A(n714), .B(n4934), .S0(n4359), .Y(n3410) );
  MXI2X1 U3783 ( .A(n713), .B(n4943), .S0(n4359), .Y(n3412) );
  MXI2X1 U3784 ( .A(n712), .B(n4913), .S0(n4359), .Y(n3414) );
  MXI2X1 U3785 ( .A(n711), .B(n4922), .S0(n4359), .Y(n3416) );
  MXI2X1 U3786 ( .A(n710), .B(n4895), .S0(n4359), .Y(n3418) );
  MXI2X1 U3787 ( .A(n709), .B(n4904), .S0(n4359), .Y(n3420) );
  MXI2X1 U3788 ( .A(n708), .B(n4874), .S0(n4359), .Y(n3422) );
  MXI2X1 U3789 ( .A(n707), .B(n4883), .S0(n4359), .Y(n3424) );
  MXI2X1 U3790 ( .A(n706), .B(n4856), .S0(n4359), .Y(n3426) );
  MXI2X1 U3791 ( .A(n705), .B(n4865), .S0(n4359), .Y(n3428) );
  MXI2X1 U3792 ( .A(n704), .B(n4834), .S0(n4360), .Y(n3430) );
  MXI2X1 U3793 ( .A(n703), .B(n4843), .S0(n4360), .Y(n3432) );
  MXI2X1 U3794 ( .A(n702), .B(n4816), .S0(n4360), .Y(n3434) );
  MXI2X1 U3795 ( .A(n701), .B(n4825), .S0(n4360), .Y(n3436) );
  MXI2X1 U3796 ( .A(n700), .B(n4790), .S0(n4360), .Y(n3438) );
  MXI2X1 U3797 ( .A(n699), .B(n4799), .S0(n4360), .Y(n3440) );
  MXI2X1 U3798 ( .A(n698), .B(n4772), .S0(n4360), .Y(n3442) );
  MXI2X1 U3799 ( .A(n697), .B(n4781), .S0(n4360), .Y(n3444) );
  MXI2X1 U3800 ( .A(n696), .B(n4750), .S0(n4360), .Y(n3446) );
  MXI2X1 U3801 ( .A(n695), .B(n4759), .S0(n4360), .Y(n3448) );
  MXI2X1 U3802 ( .A(n694), .B(n4732), .S0(n4360), .Y(n3450) );
  MXI2X1 U3803 ( .A(n693), .B(n4741), .S0(n4360), .Y(n3452) );
  MXI2X1 U3804 ( .A(n692), .B(n4710), .S0(n4359), .Y(n3454) );
  MXI2X1 U3805 ( .A(n691), .B(n4719), .S0(n4360), .Y(n3456) );
  MXI2X1 U3806 ( .A(n690), .B(n4692), .S0(n123), .Y(n3458) );
  MXI2X1 U3807 ( .A(n689), .B(n4701), .S0(n123), .Y(n3460) );
  MXI2X1 U3808 ( .A(n688), .B(n4670), .S0(n123), .Y(n3462) );
  MXI2X1 U3809 ( .A(n687), .B(n4679), .S0(n123), .Y(n3464) );
  MXI2X1 U3810 ( .A(n686), .B(n4652), .S0(n123), .Y(n3466) );
  MXI2X1 U3811 ( .A(n685), .B(n4661), .S0(n123), .Y(n3468) );
  MXI2X1 U3812 ( .A(n684), .B(n4952), .S0(n4361), .Y(n3470) );
  MXI2X1 U3813 ( .A(n683), .B(n4966), .S0(n4361), .Y(n3472) );
  MXI2X1 U3814 ( .A(n682), .B(n4934), .S0(n4361), .Y(n3474) );
  MXI2X1 U3815 ( .A(n681), .B(n4943), .S0(n4361), .Y(n3476) );
  MXI2X1 U3816 ( .A(n680), .B(n4913), .S0(n4361), .Y(n3478) );
  MXI2X1 U3817 ( .A(n679), .B(n4922), .S0(n4361), .Y(n3480) );
  MXI2X1 U3818 ( .A(n678), .B(n4895), .S0(n4361), .Y(n3482) );
  MXI2X1 U3819 ( .A(n677), .B(n4904), .S0(n4361), .Y(n3484) );
  MXI2X1 U3820 ( .A(n676), .B(n4874), .S0(n4361), .Y(n3486) );
  MXI2X1 U3821 ( .A(n675), .B(n4883), .S0(n4361), .Y(n3488) );
  MXI2X1 U3822 ( .A(n674), .B(n4856), .S0(n4361), .Y(n3490) );
  MXI2X1 U3823 ( .A(n673), .B(n4865), .S0(n4361), .Y(n3492) );
  MXI2X1 U3824 ( .A(n672), .B(n4834), .S0(n4362), .Y(n3494) );
  MXI2X1 U3825 ( .A(n671), .B(n4843), .S0(n4362), .Y(n3496) );
  MXI2X1 U3826 ( .A(n670), .B(n4816), .S0(n4362), .Y(n3498) );
  MXI2X1 U3827 ( .A(n669), .B(n4825), .S0(n4362), .Y(n3500) );
  MXI2X1 U3828 ( .A(n668), .B(n4790), .S0(n4362), .Y(n3502) );
  MXI2X1 U3829 ( .A(n667), .B(n4799), .S0(n4362), .Y(n3504) );
  MXI2X1 U3830 ( .A(n666), .B(n4772), .S0(n4362), .Y(n3506) );
  MXI2X1 U3831 ( .A(n665), .B(n4781), .S0(n4362), .Y(n3508) );
  MXI2X1 U3832 ( .A(n664), .B(n4750), .S0(n4362), .Y(n3510) );
  MXI2X1 U3833 ( .A(n663), .B(n4759), .S0(n4362), .Y(n3512) );
  MXI2X1 U3834 ( .A(n662), .B(n4732), .S0(n4362), .Y(n3514) );
  MXI2X1 U3835 ( .A(n661), .B(n4741), .S0(n4362), .Y(n3516) );
  MXI2X1 U3836 ( .A(n660), .B(n4710), .S0(n4361), .Y(n3518) );
  MXI2X1 U3837 ( .A(n659), .B(n4719), .S0(n4362), .Y(n3520) );
  MXI2X1 U3838 ( .A(n658), .B(n4692), .S0(n125), .Y(n3522) );
  MXI2X1 U3839 ( .A(n657), .B(n4701), .S0(n125), .Y(n3524) );
  MXI2X1 U3840 ( .A(n656), .B(n4670), .S0(n125), .Y(n3526) );
  MXI2X1 U3841 ( .A(n655), .B(n4679), .S0(n125), .Y(n3528) );
  MXI2X1 U3842 ( .A(n654), .B(n4652), .S0(n125), .Y(n3530) );
  MXI2X1 U3843 ( .A(n653), .B(n4661), .S0(n125), .Y(n3532) );
  CLKMX2X2 U3844 ( .A(n4570), .B(WriteData[28]), .S0(n114), .Y(n1734) );
  CLKMX2X2 U3845 ( .A(n4571), .B(WriteData[29]), .S0(n114), .Y(n1736) );
  INVXL U3846 ( .A(MEM_RegWriteData[19]), .Y(n4780) );
  INVXL U3847 ( .A(MEM_RegWriteData[17]), .Y(n4798) );
  INVXL U3848 ( .A(MEM_RegWriteData[16]), .Y(n4789) );
  INVXL U3849 ( .A(MEM_RegWriteData[18]), .Y(n4771) );
  INVXL U3850 ( .A(MEM_RegWriteData[21]), .Y(n4758) );
  INVXL U3851 ( .A(MEM_RegWriteData[20]), .Y(n4749) );
  INVXL U3852 ( .A(MEM_RegWriteData[23]), .Y(n4740) );
  INVXL U3853 ( .A(MEM_RegWriteData[22]), .Y(n4731) );
  INVXL U3854 ( .A(MEM_RegWriteData[25]), .Y(n4718) );
  INVXL U3855 ( .A(MEM_RegWriteData[24]), .Y(n4709) );
  INVXL U3856 ( .A(MEM_RegWriteData[27]), .Y(n4700) );
  INVXL U3857 ( .A(MEM_RegWriteData[26]), .Y(n4691) );
  INVXL U3858 ( .A(MEM_RegWriteData[29]), .Y(n4678) );
  INVXL U3859 ( .A(MEM_RegWriteData[28]), .Y(n4669) );
  INVXL U3860 ( .A(MEM_RegWriteData[31]), .Y(n4660) );
  INVXL U3861 ( .A(MEM_RegWriteData[30]), .Y(n4651) );
  INVXL U3862 ( .A(MEM_RegWriteData[1]), .Y(n4964) );
  INVXL U3863 ( .A(MEM_RegWriteData[0]), .Y(n4951) );
  INVXL U3864 ( .A(MEM_RegWriteData[3]), .Y(n4942) );
  INVXL U3865 ( .A(MEM_RegWriteData[2]), .Y(n4933) );
  INVXL U3866 ( .A(MEM_RegWriteData[5]), .Y(n4921) );
  INVXL U3867 ( .A(MEM_RegWriteData[4]), .Y(n4912) );
  INVXL U3868 ( .A(MEM_RegWriteData[7]), .Y(n4903) );
  INVXL U3869 ( .A(MEM_RegWriteData[6]), .Y(n4894) );
  INVXL U3870 ( .A(MEM_RegWriteData[9]), .Y(n4882) );
  INVXL U3871 ( .A(MEM_RegWriteData[8]), .Y(n4873) );
  INVXL U3872 ( .A(MEM_RegWriteData[11]), .Y(n4864) );
  INVXL U3873 ( .A(MEM_RegWriteData[10]), .Y(n4855) );
  INVXL U3874 ( .A(MEM_RegWriteData[13]), .Y(n4842) );
  INVXL U3875 ( .A(MEM_RegWriteData[12]), .Y(n4833) );
  INVXL U3876 ( .A(MEM_RegWriteData[15]), .Y(n4824) );
  INVXL U3877 ( .A(MEM_RegWriteData[14]), .Y(n4815) );
  NAND2X1 U3878 ( .A(Instruction[15]), .B(n4445), .Y(n12) );
  MXI2X1 U3879 ( .A(n4999), .B(n601), .S0(n4437), .Y(n141) );
  MXI2X1 U3880 ( .A(n4998), .B(n612), .S0(n4437), .Y(n142) );
  MXI2X1 U3881 ( .A(n4997), .B(n624), .S0(n4438), .Y(n144) );
  MXI2X1 U3882 ( .A(n4996), .B(n625), .S0(n4437), .Y(n145) );
  MXI2X1 U3883 ( .A(n4995), .B(n626), .S0(n4437), .Y(n146) );
  MXI2X1 U3884 ( .A(n4992), .B(n604), .S0(n4437), .Y(n148) );
  MXI2X1 U3885 ( .A(n4994), .B(n602), .S0(n4437), .Y(n152) );
  MXI2X1 U3886 ( .A(n4993), .B(n603), .S0(n4437), .Y(n153) );
  MXI2X1 U3887 ( .A(n4991), .B(n605), .S0(n4437), .Y(n154) );
  MXI2X1 U3888 ( .A(n4990), .B(n606), .S0(n4437), .Y(n155) );
  OAI31X1 U3889 ( .A0(n178), .A1(n179), .A2(n180), .B0(n181), .Y(n172) );
  NAND4X1 U3890 ( .A(n184), .B(n185), .C(n186), .D(n187), .Y(n178) );
  NAND4BBXL U3891 ( .AN(Instruction[15]), .BN(Instruction[26]), .C(n4998), .D(
        n183), .Y(n179) );
  NAND4X1 U3892 ( .A(n4999), .B(n4994), .C(n170), .D(n182), .Y(n180) );
  OAI22XL U3893 ( .A0(n638), .A1(n4445), .B0(n172), .B1(n4986), .Y(n3606) );
  OAI22XL U3894 ( .A0(n640), .A1(n4444), .B0(n172), .B1(n4988), .Y(n3608) );
  OAI22XL U3895 ( .A0(n641), .A1(n4444), .B0(n172), .B1(n4987), .Y(n3610) );
  NOR2BX1 U3896 ( .AN(n168), .B(n4437), .Y(n133) );
  OAI31XL U3897 ( .A0(n169), .A1(n1901), .A2(MEM_RegWrite), .B0(n167), .Y(n168) );
  OAI22XL U3898 ( .A0(n642), .A1(n4442), .B0(n176), .B1(n177), .Y(n3611) );
  NAND4X1 U3899 ( .A(n4988), .B(n4997), .C(n4996), .D(n4995), .Y(n176) );
  NAND3X1 U3900 ( .A(n4985), .B(n4986), .C(ALUOp[1]), .Y(n177) );
  CLKINVX1 U3901 ( .A(Instruction[3]), .Y(n4997) );
  CLKINVX1 U3902 ( .A(Instruction[14]), .Y(n4990) );
  CLKINVX1 U3903 ( .A(Instruction[13]), .Y(n4991) );
  CLKINVX1 U3904 ( .A(Instruction[4]), .Y(n4996) );
  CLKINVX1 U3905 ( .A(Instruction[5]), .Y(n4995) );
  CLKINVX1 U3906 ( .A(Instruction[12]), .Y(n4992) );
  CLKINVX1 U3907 ( .A(Instruction[11]), .Y(n4993) );
  CLKINVX1 U3908 ( .A(Instruction[1]), .Y(n4998) );
  CLKINVX1 U3909 ( .A(Instruction[10]), .Y(n4994) );
  CLKINVX1 U3910 ( .A(Instruction[0]), .Y(n4999) );
  OAI2BB2XL U3911 ( .B0(n639), .B1(n4445), .A0N(n4985), .A1N(ALUOp[1]), .Y(
        n3607) );
  OAI21XL U3912 ( .A0(n636), .A1(n4442), .B0(n4302), .Y(n3570) );
  OAI21XL U3913 ( .A0(n637), .A1(n4445), .B0(n4302), .Y(n3571) );
  AO22X1 U3914 ( .A0(n4441), .A1(n1939), .B0(RegDst), .B1(n4985), .Y(n3609) );
  AO22X1 U3915 ( .A0(n4640), .A1(n1), .B0(PCadd4[16]), .B1(n4363), .Y(n3572)
         );
  AO22X1 U3916 ( .A0(n4640), .A1(n2), .B0(PCadd4[17]), .B1(n4363), .Y(n3573)
         );
  AO22X1 U3917 ( .A0(n4640), .A1(n3), .B0(PCadd4[18]), .B1(n4363), .Y(n3574)
         );
  AO22X1 U3918 ( .A0(n4640), .A1(n4), .B0(PCadd4[19]), .B1(n4363), .Y(n3575)
         );
  AO22X1 U3919 ( .A0(n4640), .A1(n5), .B0(PCadd4[20]), .B1(n4363), .Y(n3576)
         );
  AO22X1 U3920 ( .A0(n4640), .A1(n6), .B0(PCadd4[21]), .B1(n4363), .Y(n3577)
         );
  AO22X1 U3921 ( .A0(n4640), .A1(n7), .B0(PCadd4[22]), .B1(n4363), .Y(n3578)
         );
  AO22X1 U3922 ( .A0(n4640), .A1(n8), .B0(PCadd4[23]), .B1(n4363), .Y(n3579)
         );
  AO22X1 U3923 ( .A0(n4364), .A1(n9), .B0(PCadd4[24]), .B1(n4363), .Y(n3580)
         );
  AO22X1 U3924 ( .A0(n4364), .A1(n11), .B0(PCadd4[25]), .B1(n4363), .Y(n3581)
         );
  AO22X1 U3925 ( .A0(n4364), .A1(n13), .B0(PCadd4[26]), .B1(n4638), .Y(n3582)
         );
  AO22X1 U3926 ( .A0(n4364), .A1(n14), .B0(PCadd4[27]), .B1(n4638), .Y(n3583)
         );
  AO22X1 U3927 ( .A0(n4364), .A1(n15), .B0(PCadd4[28]), .B1(n4638), .Y(n3584)
         );
  AO22X1 U3928 ( .A0(n4364), .A1(n16), .B0(PCadd4[29]), .B1(n4638), .Y(n3585)
         );
  AO22X1 U3929 ( .A0(n4364), .A1(n17), .B0(PCadd4[30]), .B1(n4638), .Y(n3586)
         );
  AO22X1 U3930 ( .A0(n4364), .A1(n4639), .B0(PCadd4[31]), .B1(n4638), .Y(n3587) );
  AO22X1 U3931 ( .A0(n4364), .A1(n18), .B0(PCadd4[2]), .B1(n4638), .Y(n3590)
         );
  AO22X1 U3932 ( .A0(n4364), .A1(n19), .B0(PCadd4[3]), .B1(n4638), .Y(n3591)
         );
  AO22X1 U3933 ( .A0(n4364), .A1(n20), .B0(PCadd4[4]), .B1(n4638), .Y(n3592)
         );
  AO22X1 U3934 ( .A0(n4364), .A1(n21), .B0(PCadd4[5]), .B1(n4638), .Y(n3593)
         );
  AO22X1 U3935 ( .A0(n4364), .A1(n22), .B0(PCadd4[6]), .B1(n4638), .Y(n3594)
         );
  AO22X1 U3936 ( .A0(n4364), .A1(n23), .B0(PCadd4[7]), .B1(n4638), .Y(n3595)
         );
  AO22X1 U3937 ( .A0(n4640), .A1(n24), .B0(PCadd4[8]), .B1(n4638), .Y(n3596)
         );
  AO22X1 U3938 ( .A0(n4640), .A1(n25), .B0(PCadd4[9]), .B1(n4638), .Y(n3597)
         );
  AO22X1 U3939 ( .A0(n4640), .A1(n26), .B0(PCadd4[10]), .B1(n4638), .Y(n3598)
         );
  AO22X1 U3940 ( .A0(n4640), .A1(n27), .B0(PCadd4[11]), .B1(n4638), .Y(n3599)
         );
  AO22X1 U3941 ( .A0(n4640), .A1(n28), .B0(PCadd4[12]), .B1(n4363), .Y(n3600)
         );
  AO22X1 U3942 ( .A0(n4640), .A1(n29), .B0(PCadd4[13]), .B1(n4363), .Y(n3601)
         );
  AO22X1 U3943 ( .A0(n4640), .A1(n30), .B0(PCadd4[14]), .B1(n4363), .Y(n3602)
         );
  AO22X1 U3944 ( .A0(n4640), .A1(n31), .B0(PCadd4[15]), .B1(n4363), .Y(n3603)
         );
  AO22X1 U3945 ( .A0(n4441), .A1(EX[0]), .B0(ALUSrc), .B1(n4985), .Y(n3605) );
  AO22X1 U3946 ( .A0(n4441), .A1(MEM[0]), .B0(MemWrite), .B1(n4985), .Y(n3612)
         );
  AO22X1 U3947 ( .A0(n4441), .A1(MEM[1]), .B0(MemRead), .B1(n4985), .Y(n3613)
         );
  AO22X1 U3948 ( .A0(n4441), .A1(WB[0]), .B0(MemtoReg), .B1(n4985), .Y(n3614)
         );
  AO22X1 U3949 ( .A0(n4441), .A1(WB[1]), .B0(RegWrite), .B1(n4985), .Y(n3615)
         );
  AO22X1 U3950 ( .A0(n4640), .A1(n32), .B0(PCadd4[0]), .B1(n4638), .Y(n3588)
         );
  AO22X1 U3951 ( .A0(n4640), .A1(n33), .B0(PCadd4[1]), .B1(n4638), .Y(n3589)
         );
  NOR4X1 U3952 ( .A(Instruction[14]), .B(Instruction[13]), .C(Instruction[12]), 
        .D(Instruction[11]), .Y(n182) );
  OAI22XL U3953 ( .A0(n633), .A1(n4445), .B0(n4437), .B1(n4991), .Y(n3567) );
  OAI22XL U3954 ( .A0(n634), .A1(n4443), .B0(n4436), .B1(n4990), .Y(n3568) );
  OAI22XL U3955 ( .A0(n631), .A1(n4445), .B0(n4437), .B1(n4993), .Y(n3565) );
  OAI22XL U3956 ( .A0(n632), .A1(n4446), .B0(n4436), .B1(n4992), .Y(n3566) );
  NOR3X1 U3957 ( .A(Instruction[5]), .B(Instruction[7]), .C(Instruction[6]), 
        .Y(n184) );
  MXI2X1 U3958 ( .A(n4423), .B(n643), .S0(n4436), .Y(n3616) );
  MXI2X1 U3959 ( .A(n4424), .B(n644), .S0(n4436), .Y(n3617) );
  MXI2X1 U3960 ( .A(n4425), .B(n645), .S0(n4436), .Y(n3618) );
  MXI2X1 U3961 ( .A(n4427), .B(n646), .S0(n4436), .Y(n3619) );
  MXI2X1 U3962 ( .A(n4428), .B(n647), .S0(n4436), .Y(n3620) );
  MXI2X1 U3963 ( .A(n4430), .B(n648), .S0(n4436), .Y(n3621) );
  MXI2X1 U3964 ( .A(n4431), .B(n649), .S0(n4436), .Y(n3622) );
  MXI2X1 U3965 ( .A(n4432), .B(n650), .S0(n4436), .Y(n3623) );
  MXI2X1 U3966 ( .A(n4434), .B(n651), .S0(n4436), .Y(n3624) );
  MXI2X1 U3967 ( .A(n4435), .B(n652), .S0(n4436), .Y(n3625) );
  OAI21XL U3968 ( .A0(n1899), .A1(n133), .B0(n134), .Y(n3604) );
  OAI21XL U3969 ( .A0(n635), .A1(n4447), .B0(n12), .Y(n3569) );
  CLKINVX3 U3970 ( .A(WriteData[0]), .Y(n4952) );
  CLKINVX3 U3971 ( .A(WriteData[1]), .Y(n4966) );
  CLKINVX3 U3972 ( .A(WriteData[2]), .Y(n4934) );
  CLKINVX3 U3973 ( .A(WriteData[3]), .Y(n4943) );
  CLKINVX3 U3974 ( .A(WriteData[4]), .Y(n4913) );
  CLKINVX3 U3975 ( .A(WriteData[5]), .Y(n4922) );
  CLKINVX3 U3976 ( .A(WriteData[6]), .Y(n4895) );
  CLKINVX3 U3977 ( .A(WriteData[7]), .Y(n4904) );
  CLKINVX3 U3978 ( .A(WriteData[8]), .Y(n4874) );
  CLKINVX3 U3979 ( .A(WriteData[9]), .Y(n4883) );
  CLKINVX3 U3980 ( .A(WriteData[10]), .Y(n4856) );
  CLKINVX3 U3981 ( .A(WriteData[11]), .Y(n4865) );
  CLKINVX3 U3982 ( .A(WriteData[12]), .Y(n4834) );
  CLKINVX3 U3983 ( .A(WriteData[13]), .Y(n4843) );
  CLKINVX3 U3984 ( .A(WriteData[14]), .Y(n4816) );
  CLKINVX3 U3985 ( .A(WriteData[15]), .Y(n4825) );
  CLKINVX3 U3986 ( .A(WriteData[16]), .Y(n4790) );
  CLKINVX3 U3987 ( .A(WriteData[17]), .Y(n4799) );
  CLKINVX3 U3988 ( .A(WriteData[18]), .Y(n4772) );
  CLKINVX3 U3989 ( .A(WriteData[19]), .Y(n4781) );
  CLKINVX3 U3990 ( .A(WriteData[20]), .Y(n4750) );
  CLKINVX3 U3991 ( .A(WriteData[21]), .Y(n4759) );
  CLKINVX3 U3992 ( .A(WriteData[22]), .Y(n4732) );
  CLKINVX3 U3993 ( .A(WriteData[23]), .Y(n4741) );
  CLKINVX3 U3994 ( .A(WriteData[24]), .Y(n4710) );
  CLKINVX3 U3995 ( .A(WriteData[25]), .Y(n4719) );
  CLKINVX3 U3996 ( .A(WriteData[26]), .Y(n4692) );
  CLKINVX3 U3997 ( .A(WriteData[27]), .Y(n4701) );
  CLKINVX3 U3998 ( .A(WriteData[28]), .Y(n4670) );
  CLKINVX3 U3999 ( .A(WriteData[29]), .Y(n4679) );
  CLKINVX3 U4000 ( .A(WriteData[30]), .Y(n4652) );
  CLKINVX3 U4001 ( .A(WriteData[31]), .Y(n4661) );
  CLKINVX3 U4002 ( .A(n124), .Y(n4574) );
  CLKINVX3 U4003 ( .A(n133), .Y(n4640) );
  CLKINVX3 U4004 ( .A(n134), .Y(n4638) );
  InstructionDecode_DW_mult_uns_1 mult_add_145_aco ( .a({
        next_Immediate_SE[29:15], n155, n154, n148, n153, n152, n151, n147, 
        n150, n149, n146, n145, n144, n143, n142, n141, 1'b0, 1'b0}), .b(n1795), .product({SYNOPSYS_UNCONNECTED__0, N484, N483, N482, N481, N480, N479, N478, 
        N477, N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, 
        N465, N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2}) );
  InstructionDecode_DW01_add_2 add_145_aco ( .A(PCadd4), .B({N484, N483, N482, 
        N481, N480, N479, N478, N477, N476, N475, N474, N473, N472, N471, N470, 
        N469, N468, N467, N466, N465, N464, N463, N462, N461, N460, N459, N458, 
        N457, N456, N455, 1'b0, 1'b0}), .CI(1'b0), .SUM(PCbranched) );
  SDFFRXL \EX_reg[6]  ( .D(n3611), .SI(EX[5]), .SE(test_se), .CK(clk), .RN(
        n4451), .Q(EX[6]), .QN(n642) );
  SDFFRXL \EX_reg[5]  ( .D(n3610), .SI(n37), .SE(test_se), .CK(clk), .RN(n4451), .Q(EX[5]), .QN(n641) );
  SDFFRXL \WB_reg[0]  ( .D(n3614), .SI(n647), .SE(test_se), .CK(clk), .RN(
        n4450), .Q(WB[0]), .QN(n1753) );
  SDFFRXL \MEM_reg[0]  ( .D(n3612), .SI(n637), .SE(test_se), .CK(clk), .RN(
        n4451), .Q(MEM[0]), .QN(n1751) );
  SDFFRXL \WB_reg[1]  ( .D(n3615), .SI(n1753), .SE(test_se), .CK(clk), .RN(
        n4450), .Q(WB[1]), .QN(test_so2) );
  SDFFRXL \RegisterRd_reg[4]  ( .D(n3569), .SI(n634), .SE(test_se), .CK(clk), 
        .RN(n4462), .Q(RegisterRd[4]), .QN(n635) );
  SDFFRXL \RegisterRd_reg[1]  ( .D(n3566), .SI(n631), .SE(test_se), .CK(clk), 
        .RN(n4462), .Q(RegisterRd[1]), .QN(n632) );
  SDFFRXL \RegisterRd_reg[3]  ( .D(n3568), .SI(n633), .SE(test_se), .CK(clk), 
        .RN(n4462), .Q(RegisterRd[3]), .QN(n634) );
  SDFFRXL \RegisterRd_reg[2]  ( .D(n3567), .SI(n632), .SE(test_se), .CK(clk), 
        .RN(n4462), .Q(RegisterRd[2]), .QN(n633) );
  SDFFRXL \RegisterRd_reg[0]  ( .D(n3565), .SI(n67), .SE(test_se), .CK(clk), 
        .RN(n4462), .Q(RegisterRd[0]), .QN(n631) );
  SDFFRXL \Immediate_SE_reg[31]  ( .D(n3571), .SI(n636), .SE(test_se), .CK(clk), .RN(n4459), .Q(Immediate_SE[31]), .QN(n637) );
  SDFFRXL \Immediate_SE_reg[30]  ( .D(n3570), .SI(n622), .SE(test_se), .CK(clk), .RN(n4459), .Q(Immediate_SE[30]), .QN(n636) );
  SDFFRXL \Immediate_SE_reg[29]  ( .D(next_Immediate_SE[29]), .SI(n621), .SE(
        test_se), .CK(clk), .RN(n4460), .Q(Immediate_SE[29]), .QN(n622) );
  SDFFRXL \Immediate_SE_reg[28]  ( .D(next_Immediate_SE[28]), .SI(n620), .SE(
        test_se), .CK(clk), .RN(n4460), .Q(Immediate_SE[28]), .QN(n621) );
  SDFFRXL \Immediate_SE_reg[27]  ( .D(next_Immediate_SE[27]), .SI(n619), .SE(
        test_se), .CK(clk), .RN(n4460), .Q(Immediate_SE[27]), .QN(n620) );
  SDFFRXL \Immediate_SE_reg[26]  ( .D(next_Immediate_SE[26]), .SI(n618), .SE(
        test_se), .CK(clk), .RN(n4460), .Q(Immediate_SE[26]), .QN(n619) );
  SDFFRXL \Immediate_SE_reg[23]  ( .D(next_Immediate_SE[23]), .SI(n615), .SE(
        test_se), .CK(clk), .RN(n4460), .Q(Immediate_SE[23]), .QN(n616) );
  SDFFRXL \Immediate_SE_reg[22]  ( .D(next_Immediate_SE[22]), .SI(n614), .SE(
        test_se), .CK(clk), .RN(n4460), .Q(Immediate_SE[22]), .QN(n615) );
  SDFFRXL \Immediate_SE_reg[21]  ( .D(next_Immediate_SE[21]), .SI(n613), .SE(
        test_se), .CK(clk), .RN(n4460), .Q(Immediate_SE[21]), .QN(n614) );
  SDFFRXL \Immediate_SE_reg[19]  ( .D(next_Immediate_SE[19]), .SI(n610), .SE(
        test_se), .CK(clk), .RN(n4460), .Q(Immediate_SE[19]), .QN(n611) );
  SDFFRXL \Immediate_SE_reg[18]  ( .D(next_Immediate_SE[18]), .SI(n609), .SE(
        test_se), .CK(clk), .RN(n4460), .Q(Immediate_SE[18]), .QN(n610) );
  SDFFRXL \Immediate_SE_reg[17]  ( .D(next_Immediate_SE[17]), .SI(n608), .SE(
        test_se), .CK(clk), .RN(n4461), .Q(Immediate_SE[17]), .QN(n609) );
  SDFFRXL \Immediate_SE_reg[16]  ( .D(next_Immediate_SE[16]), .SI(n607), .SE(
        test_se), .CK(clk), .RN(n4461), .Q(Immediate_SE[16]), .QN(n608) );
  SDFFRXL \Immediate_SE_reg[12]  ( .D(n148), .SI(n603), .SE(test_se), .CK(clk), 
        .RN(n4461), .Q(Immediate_SE[12]), .QN(n604) );
  SDFFRXL \EX_reg[3]  ( .D(n3608), .SI(n639), .SE(test_se), .CK(clk), .RN(
        n4451), .Q(EX[3]), .QN(n640) );
  SDFFRXL \PCBuffer_reg[15]  ( .D(n3603), .SI(n30), .SE(test_se), .CK(clk), 
        .RN(n4451), .Q(n31), .QN(n3642) );
  SDFFRXL \PCBuffer_reg[14]  ( .D(n3602), .SI(n29), .SE(test_se), .CK(clk), 
        .RN(n4451), .Q(n30), .QN(n3643) );
  SDFFRXL \PCBuffer_reg[13]  ( .D(n3601), .SI(n28), .SE(test_se), .CK(clk), 
        .RN(n4452), .Q(n29), .QN(n3644) );
  SDFFRXL \PCBuffer_reg[12]  ( .D(n3600), .SI(n27), .SE(test_se), .CK(clk), 
        .RN(n4452), .Q(n28), .QN(n3645) );
  SDFFRXL \PCBuffer_reg[11]  ( .D(n3599), .SI(n26), .SE(test_se), .CK(clk), 
        .RN(n4452), .Q(n27), .QN(n3646) );
  SDFFRXL \PCBuffer_reg[10]  ( .D(n3598), .SI(n25), .SE(test_se), .CK(clk), 
        .RN(n4452), .Q(n26), .QN(n3647) );
  SDFFRXL \PCBuffer_reg[9]  ( .D(n3597), .SI(n24), .SE(test_se), .CK(clk), 
        .RN(n4452), .Q(n25), .QN(n3648) );
  SDFFRXL \PCBuffer_reg[8]  ( .D(n3596), .SI(n23), .SE(test_se), .CK(clk), 
        .RN(n4452), .Q(n24), .QN(n3649) );
  SDFFRXL \PCBuffer_reg[7]  ( .D(n3595), .SI(n22), .SE(test_se), .CK(clk), 
        .RN(n4452), .Q(n23), .QN(n3650) );
  SDFFRXL \PCBuffer_reg[6]  ( .D(n3594), .SI(n21), .SE(test_se), .CK(clk), 
        .RN(n4452), .Q(n22), .QN(n3651) );
  SDFFRXL \PCBuffer_reg[5]  ( .D(n3593), .SI(n20), .SE(test_se), .CK(clk), 
        .RN(n4452), .Q(n21), .QN(n3652) );
  SDFFRXL \PCBuffer_reg[4]  ( .D(n3592), .SI(n19), .SE(test_se), .CK(clk), 
        .RN(n4452), .Q(n20), .QN(n3653) );
  SDFFRXL \PCBuffer_reg[3]  ( .D(n3591), .SI(n18), .SE(test_se), .CK(clk), 
        .RN(n4452), .Q(n19), .QN(n3654) );
  SDFFRXL \PCBuffer_reg[2]  ( .D(n3590), .SI(n33), .SE(test_se), .CK(clk), 
        .RN(n4452), .Q(n18), .QN(n3655) );
  SDFFRXL \PCBuffer_reg[1]  ( .D(n3589), .SI(n32), .SE(test_se), .CK(clk), 
        .RN(n4453), .Q(n33), .QN(n3656) );
  SDFFRXL \PCBuffer_reg[0]  ( .D(n3588), .SI(n1743), .SE(test_se), .CK(clk), 
        .RN(n4453), .Q(n32), .QN(n3657) );
  SDFFRXL \PCBuffer_reg[30]  ( .D(n3586), .SI(n16), .SE(test_se), .CK(clk), 
        .RN(n4453), .Q(n17), .QN(n3627) );
  SDFFRXL \PCBuffer_reg[29]  ( .D(n3585), .SI(n15), .SE(test_se), .CK(clk), 
        .RN(n4453), .Q(n16), .QN(n3628) );
  SDFFRXL \PCBuffer_reg[28]  ( .D(n3584), .SI(n14), .SE(test_se), .CK(clk), 
        .RN(n4453), .Q(n15), .QN(n3629) );
  SDFFRXL \PCBuffer_reg[27]  ( .D(n3583), .SI(n13), .SE(test_se), .CK(clk), 
        .RN(n4453), .Q(n14), .QN(n3630) );
  SDFFRXL \PCBuffer_reg[26]  ( .D(n3582), .SI(n11), .SE(test_se), .CK(clk), 
        .RN(n4453), .Q(n13), .QN(n3631) );
  SDFFRXL \PCBuffer_reg[25]  ( .D(n3581), .SI(n9), .SE(test_se), .CK(clk), 
        .RN(n4453), .Q(n11), .QN(n3632) );
  SDFFRXL \PCBuffer_reg[24]  ( .D(n3580), .SI(n8), .SE(test_se), .CK(clk), 
        .RN(n4453), .Q(n9), .QN(n3633) );
  SDFFRXL \PCBuffer_reg[23]  ( .D(n3579), .SI(n7), .SE(test_se), .CK(clk), 
        .RN(n4453), .Q(n8), .QN(n3634) );
  SDFFRXL \PCBuffer_reg[22]  ( .D(n3578), .SI(n6), .SE(test_se), .CK(clk), 
        .RN(n4453), .Q(n7), .QN(n3635) );
  SDFFRXL \PCBuffer_reg[21]  ( .D(n3577), .SI(n5), .SE(test_se), .CK(clk), 
        .RN(n4454), .Q(n6), .QN(n3636) );
  SDFFRXL \PCBuffer_reg[20]  ( .D(n3576), .SI(n4), .SE(test_se), .CK(clk), 
        .RN(n4454), .Q(n5), .QN(n3637) );
  SDFFRXL \PCBuffer_reg[19]  ( .D(n3575), .SI(n3), .SE(test_se), .CK(clk), 
        .RN(n4454), .Q(n4), .QN(n3638) );
  SDFFRXL \PCBuffer_reg[18]  ( .D(n3574), .SI(n2), .SE(test_se), .CK(clk), 
        .RN(n4454), .Q(n3), .QN(n3639) );
  SDFFRXL \PCBuffer_reg[17]  ( .D(n3573), .SI(n1), .SE(test_se), .CK(clk), 
        .RN(n4454), .Q(n2), .QN(n3640) );
  SDFFRXL \PCBuffer_reg[16]  ( .D(n3572), .SI(n31), .SE(test_se), .CK(clk), 
        .RN(n4454), .Q(n1), .QN(n3641) );
  SDFFRXL \MEM_reg[1]  ( .D(n3613), .SI(n1751), .SE(test_se), .CK(clk), .RN(
        n4451), .Q(MEM[1]), .QN(n1743) );
  SDFFRXL \Immediate_SE_reg[0]  ( .D(n141), .SI(EX[6]), .SE(test_se), .CK(clk), 
        .RN(n4462), .Q(Immediate_SE[0]), .QN(n601) );
  SDFFRXL \EX_reg[1]  ( .D(n3606), .SI(n38), .SE(test_se), .CK(clk), .RN(n4451), .Q(n1945), .QN(n638) );
  SDFFRXL \Immediate_SE_reg[15]  ( .D(next_Immediate_SE[15]), .SI(n606), .SE(
        test_se), .CK(clk), .RN(n4461), .Q(Immediate_SE[15]), .QN(n607) );
  SDFFRXL \Immediate_SE_reg[14]  ( .D(n155), .SI(n605), .SE(test_se), .CK(clk), 
        .RN(n4461), .Q(Immediate_SE[14]), .QN(n606) );
  SDFFRXL \Immediate_SE_reg[13]  ( .D(n154), .SI(n604), .SE(test_se), .CK(clk), 
        .RN(n4461), .Q(Immediate_SE[13]), .QN(n605) );
  SDFFRXL \Immediate_SE_reg[11]  ( .D(n153), .SI(n602), .SE(test_se), .CK(clk), 
        .RN(n4461), .Q(Immediate_SE[11]), .QN(n603) );
  SDFFRXL \Immediate_SE_reg[10]  ( .D(n152), .SI(n1675), .SE(test_se), .CK(clk), .RN(n4461), .Q(Immediate_SE[10]), .QN(n602) );
  SDFFRXL \Immediate_SE_reg[9]  ( .D(n151), .SI(n1673), .SE(test_se), .CK(clk), 
        .RN(n4461), .Q(Immediate_SE[9]), .QN(n1675) );
  SDFFRXL \Immediate_SE_reg[8]  ( .D(n147), .SI(n1671), .SE(test_se), .CK(clk), 
        .RN(n4461), .Q(Immediate_SE[8]), .QN(n1673) );
  SDFFRXL \Immediate_SE_reg[7]  ( .D(n150), .SI(n1669), .SE(test_se), .CK(clk), 
        .RN(n4461), .Q(Immediate_SE[7]), .QN(n1671) );
  SDFFRXL \Immediate_SE_reg[6]  ( .D(n149), .SI(n626), .SE(test_se), .CK(clk), 
        .RN(n4461), .Q(Immediate_SE[6]), .QN(n1669) );
  SDFFRXL \Immediate_SE_reg[4]  ( .D(n145), .SI(n624), .SE(test_se), .CK(clk), 
        .RN(n4462), .Q(Immediate_SE[4]), .QN(n625) );
  SDFFRXL PCBuffer_valid_reg ( .D(n3604), .SI(n4639), .SE(test_se), .CK(clk), 
        .RN(n4451), .Q(PCBuffer_valid), .QN(n3658) );
  SDFFRXL \Immediate_SE_reg[3]  ( .D(n144), .SI(n39), .SE(test_se), .CK(clk), 
        .RN(n4462), .Q(Immediate_SE[3]), .QN(n624) );
  SDFFRXL \RegisterRs_reg[4]  ( .D(n3625), .SI(n651), .SE(test_se), .CK(clk), 
        .RN(n4450), .Q(RegisterRs[4]), .QN(n652) );
  SDFFNSRXL \regfile_reg[31][31]  ( .D(n3690), .SI(n570), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4462), .Q(\regfile[31][31] ), .QN(n569) );
  SDFFNSRXL \regfile_reg[31][30]  ( .D(n3689), .SI(n571), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4462), .Q(\regfile[31][30] ), .QN(n570) );
  SDFFNSRXL \regfile_reg[31][29]  ( .D(n3688), .SI(n572), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4463), .Q(\regfile[31][29] ), .QN(n571) );
  SDFFNSRXL \regfile_reg[31][28]  ( .D(n3687), .SI(n573), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4463), .Q(\regfile[31][28] ), .QN(n572) );
  SDFFNSRXL \regfile_reg[31][27]  ( .D(n3686), .SI(n574), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4463), .Q(\regfile[31][27] ), .QN(n573) );
  SDFFNSRXL \regfile_reg[31][26]  ( .D(n3685), .SI(n575), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4463), .Q(\regfile[31][26] ), .QN(n574) );
  SDFFNSRXL \regfile_reg[31][25]  ( .D(n3684), .SI(n576), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4463), .Q(\regfile[31][25] ), .QN(n575) );
  SDFFNSRXL \regfile_reg[31][24]  ( .D(n3683), .SI(n577), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4463), .Q(\regfile[31][24] ), .QN(n576) );
  SDFFNSRXL \regfile_reg[31][23]  ( .D(n3682), .SI(n578), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4463), .Q(\regfile[31][23] ), .QN(n577) );
  SDFFNSRXL \regfile_reg[31][22]  ( .D(n3681), .SI(n579), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4463), .Q(\regfile[31][22] ), .QN(n578) );
  SDFFNSRXL \regfile_reg[31][21]  ( .D(n3680), .SI(n580), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4463), .Q(\regfile[31][21] ), .QN(n579) );
  SDFFNSRXL \regfile_reg[31][20]  ( .D(n3679), .SI(n581), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4463), .Q(\regfile[31][20] ), .QN(n580) );
  SDFFNSRXL \regfile_reg[31][19]  ( .D(n3678), .SI(n582), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4463), .Q(\regfile[31][19] ), .QN(n581) );
  SDFFNSRXL \regfile_reg[31][18]  ( .D(n3677), .SI(n583), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4463), .Q(\regfile[31][18] ), .QN(n582) );
  SDFFNSRXL \regfile_reg[31][17]  ( .D(n3676), .SI(n584), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4463), .Q(\regfile[31][17] ), .QN(n583) );
  SDFFNSRXL \regfile_reg[31][16]  ( .D(n3675), .SI(n585), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4463), .Q(\regfile[31][16] ), .QN(n584) );
  SDFFNSRXL \regfile_reg[31][15]  ( .D(n3674), .SI(n586), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4463), .Q(\regfile[31][15] ), .QN(n585) );
  SDFFNSRXL \regfile_reg[31][14]  ( .D(n3673), .SI(n587), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4463), .Q(\regfile[31][14] ), .QN(n586) );
  SDFFNSRXL \regfile_reg[31][13]  ( .D(n3672), .SI(n588), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4463), .Q(\regfile[31][13] ), .QN(n587) );
  SDFFNSRXL \regfile_reg[31][12]  ( .D(n3671), .SI(n589), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4463), .Q(\regfile[31][12] ), .QN(n588) );
  SDFFNSRXL \regfile_reg[31][11]  ( .D(n3670), .SI(n590), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4464), .Q(\regfile[31][11] ), .QN(n589) );
  SDFFNSRXL \regfile_reg[31][10]  ( .D(n3669), .SI(n591), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4464), .Q(\regfile[31][10] ), .QN(n590) );
  SDFFNSRXL \regfile_reg[31][9]  ( .D(n3668), .SI(n592), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4464), .Q(\regfile[31][9] ), .QN(n591) );
  SDFFNSRXL \regfile_reg[31][8]  ( .D(n3667), .SI(n593), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4464), .Q(\regfile[31][8] ), .QN(n592) );
  SDFFNSRXL \regfile_reg[31][7]  ( .D(n3666), .SI(n594), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4464), .Q(\regfile[31][7] ), .QN(n593) );
  SDFFNSRXL \regfile_reg[31][6]  ( .D(n3665), .SI(n595), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4464), .Q(\regfile[31][6] ), .QN(n594) );
  SDFFNSRXL \regfile_reg[31][5]  ( .D(n3664), .SI(n596), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4464), .Q(\regfile[31][5] ), .QN(n595) );
  SDFFNSRXL \regfile_reg[31][4]  ( .D(n3663), .SI(n597), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4464), .Q(\regfile[31][4] ), .QN(n596) );
  SDFFNSRXL \regfile_reg[31][3]  ( .D(n3662), .SI(n598), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4464), .Q(\regfile[31][3] ), .QN(n597) );
  SDFFNSRXL \regfile_reg[31][2]  ( .D(n3661), .SI(n599), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4464), .Q(\regfile[31][2] ), .QN(n598) );
  SDFFNSRXL \regfile_reg[31][1]  ( .D(n3660), .SI(n600), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4464), .Q(\regfile[31][1] ), .QN(n599) );
  SDFFNSRXL \regfile_reg[31][0]  ( .D(n3659), .SI(n653), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4464), .Q(\regfile[31][0] ), .QN(n600) );
  SDFFNSRXL \regfile_reg[27][31]  ( .D(n3340), .SI(n750), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4470), .Q(\regfile[27][31] ), .QN(n749) );
  SDFFNSRXL \regfile_reg[27][30]  ( .D(n3338), .SI(n751), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4470), .Q(\regfile[27][30] ), .QN(n750) );
  SDFFNSRXL \regfile_reg[27][29]  ( .D(n3336), .SI(n752), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4470), .Q(\regfile[27][29] ), .QN(n751) );
  SDFFNSRXL \regfile_reg[27][28]  ( .D(n3334), .SI(n753), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4470), .Q(\regfile[27][28] ), .QN(n752) );
  SDFFNSRXL \regfile_reg[27][27]  ( .D(n3332), .SI(n754), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4470), .Q(\regfile[27][27] ), .QN(n753) );
  SDFFNSRXL \regfile_reg[27][26]  ( .D(n3330), .SI(n755), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4470), .Q(\regfile[27][26] ), .QN(n754) );
  SDFFNSRXL \regfile_reg[27][25]  ( .D(n3328), .SI(n756), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4470), .Q(\regfile[27][25] ), .QN(n755) );
  SDFFNSRXL \regfile_reg[27][24]  ( .D(n3326), .SI(n757), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4470), .Q(\regfile[27][24] ), .QN(n756) );
  SDFFNSRXL \regfile_reg[27][23]  ( .D(n3324), .SI(n758), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4470), .Q(\regfile[27][23] ), .QN(n757) );
  SDFFNSRXL \regfile_reg[27][22]  ( .D(n3322), .SI(n759), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4470), .Q(\regfile[27][22] ), .QN(n758) );
  SDFFNSRXL \regfile_reg[27][21]  ( .D(n3320), .SI(n760), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4470), .Q(\regfile[27][21] ), .QN(n759) );
  SDFFNSRXL \regfile_reg[27][20]  ( .D(n3318), .SI(n761), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4470), .Q(\regfile[27][20] ), .QN(n760) );
  SDFFNSRXL \regfile_reg[27][19]  ( .D(n3316), .SI(n762), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4470), .Q(\regfile[27][19] ), .QN(n761) );
  SDFFNSRXL \regfile_reg[27][18]  ( .D(n3314), .SI(n763), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4470), .Q(\regfile[27][18] ), .QN(n762) );
  SDFFNSRXL \regfile_reg[27][17]  ( .D(n3312), .SI(n764), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4470), .Q(\regfile[27][17] ), .QN(n763) );
  SDFFNSRXL \regfile_reg[27][16]  ( .D(n3310), .SI(n765), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4470), .Q(\regfile[27][16] ), .QN(n764) );
  SDFFNSRXL \regfile_reg[27][15]  ( .D(n3308), .SI(n766), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4470), .Q(\regfile[27][15] ), .QN(n765) );
  SDFFNSRXL \regfile_reg[27][14]  ( .D(n3306), .SI(n767), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4470), .Q(\regfile[27][14] ), .QN(n766) );
  SDFFNSRXL \regfile_reg[27][13]  ( .D(n3304), .SI(n768), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4471), .Q(\regfile[27][13] ), .QN(n767) );
  SDFFNSRXL \regfile_reg[27][12]  ( .D(n3302), .SI(n769), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4471), .Q(\regfile[27][12] ), .QN(n768) );
  SDFFNSRXL \regfile_reg[27][11]  ( .D(n3300), .SI(n770), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4471), .Q(\regfile[27][11] ), .QN(n769) );
  SDFFNSRXL \regfile_reg[27][10]  ( .D(n3298), .SI(n771), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4471), .Q(\regfile[27][10] ), .QN(n770) );
  SDFFNSRXL \regfile_reg[27][9]  ( .D(n3296), .SI(n772), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4471), .Q(\regfile[27][9] ), .QN(n771) );
  SDFFNSRXL \regfile_reg[27][8]  ( .D(n3294), .SI(n773), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4471), .Q(\regfile[27][8] ), .QN(n772) );
  SDFFNSRXL \regfile_reg[27][7]  ( .D(n3292), .SI(n774), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4471), .Q(\regfile[27][7] ), .QN(n773) );
  SDFFNSRXL \regfile_reg[27][6]  ( .D(n3290), .SI(n775), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4471), .Q(\regfile[27][6] ), .QN(n774) );
  SDFFNSRXL \regfile_reg[27][5]  ( .D(n3288), .SI(n776), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4471), .Q(\regfile[27][5] ), .QN(n775) );
  SDFFNSRXL \regfile_reg[27][4]  ( .D(n3286), .SI(n777), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4471), .Q(\regfile[27][4] ), .QN(n776) );
  SDFFNSRXL \regfile_reg[27][3]  ( .D(n3284), .SI(n778), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4471), .Q(\regfile[27][3] ), .QN(n777) );
  SDFFNSRXL \regfile_reg[27][2]  ( .D(n3282), .SI(n779), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4471), .Q(\regfile[27][2] ), .QN(n778) );
  SDFFNSRXL \regfile_reg[27][1]  ( .D(n3280), .SI(n780), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4471), .Q(\regfile[27][1] ), .QN(n779) );
  SDFFNSRXL \regfile_reg[27][0]  ( .D(n3278), .SI(n781), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4471), .Q(\regfile[27][0] ), .QN(n780) );
  SDFFNSRXL \regfile_reg[23][31]  ( .D(n3084), .SI(n878), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4477), .Q(\regfile[23][31] ), .QN(n877) );
  SDFFNSRXL \regfile_reg[23][30]  ( .D(n3082), .SI(n879), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4477), .Q(\regfile[23][30] ), .QN(n878) );
  SDFFNSRXL \regfile_reg[23][29]  ( .D(n3080), .SI(n880), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4477), .Q(\regfile[23][29] ), .QN(n879) );
  SDFFNSRXL \regfile_reg[23][28]  ( .D(n3078), .SI(n881), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4477), .Q(\regfile[23][28] ), .QN(n880) );
  SDFFNSRXL \regfile_reg[23][27]  ( .D(n3076), .SI(n882), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4477), .Q(\regfile[23][27] ), .QN(n881) );
  SDFFNSRXL \regfile_reg[23][26]  ( .D(n3074), .SI(n883), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4477), .Q(\regfile[23][26] ), .QN(n882) );
  SDFFNSRXL \regfile_reg[23][25]  ( .D(n3072), .SI(n884), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4477), .Q(\regfile[23][25] ), .QN(n883) );
  SDFFNSRXL \regfile_reg[23][24]  ( .D(n3070), .SI(n885), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4477), .Q(\regfile[23][24] ), .QN(n884) );
  SDFFNSRXL \regfile_reg[23][23]  ( .D(n3068), .SI(n886), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4477), .Q(\regfile[23][23] ), .QN(n885) );
  SDFFNSRXL \regfile_reg[23][22]  ( .D(n3066), .SI(n887), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4477), .Q(\regfile[23][22] ), .QN(n886) );
  SDFFNSRXL \regfile_reg[23][21]  ( .D(n3064), .SI(n888), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4477), .Q(\regfile[23][21] ), .QN(n887) );
  SDFFNSRXL \regfile_reg[23][20]  ( .D(n3062), .SI(n889), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4477), .Q(\regfile[23][20] ), .QN(n888) );
  SDFFNSRXL \regfile_reg[23][19]  ( .D(n3060), .SI(n890), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4477), .Q(\regfile[23][19] ), .QN(n889) );
  SDFFNSRXL \regfile_reg[23][18]  ( .D(n3058), .SI(n891), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4477), .Q(\regfile[23][18] ), .QN(n890) );
  SDFFNSRXL \regfile_reg[23][17]  ( .D(n3056), .SI(n892), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4477), .Q(\regfile[23][17] ), .QN(n891) );
  SDFFNSRXL \regfile_reg[23][16]  ( .D(n3054), .SI(n893), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4477), .Q(\regfile[23][16] ), .QN(n892) );
  SDFFNSRXL \regfile_reg[23][15]  ( .D(n3052), .SI(n894), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4478), .Q(\regfile[23][15] ), .QN(n893) );
  SDFFNSRXL \regfile_reg[23][14]  ( .D(n3050), .SI(n895), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4478), .Q(\regfile[23][14] ), .QN(n894) );
  SDFFNSRXL \regfile_reg[23][13]  ( .D(n3048), .SI(n896), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4478), .Q(\regfile[23][13] ), .QN(n895) );
  SDFFNSRXL \regfile_reg[23][12]  ( .D(n3046), .SI(n897), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4478), .Q(\regfile[23][12] ), .QN(n896) );
  SDFFNSRXL \regfile_reg[23][11]  ( .D(n3044), .SI(n898), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4478), .Q(\regfile[23][11] ), .QN(n897) );
  SDFFNSRXL \regfile_reg[23][10]  ( .D(n3042), .SI(n899), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4478), .Q(\regfile[23][10] ), .QN(n898) );
  SDFFNSRXL \regfile_reg[23][9]  ( .D(n3040), .SI(n900), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4478), .Q(\regfile[23][9] ), .QN(n899) );
  SDFFNSRXL \regfile_reg[23][8]  ( .D(n3038), .SI(n901), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4478), .Q(\regfile[23][8] ), .QN(n900) );
  SDFFNSRXL \regfile_reg[23][7]  ( .D(n3036), .SI(n902), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4478), .Q(\regfile[23][7] ), .QN(n901) );
  SDFFNSRXL \regfile_reg[23][6]  ( .D(n3034), .SI(n903), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4478), .Q(\regfile[23][6] ), .QN(n902) );
  SDFFNSRXL \regfile_reg[23][5]  ( .D(n3032), .SI(n904), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4478), .Q(\regfile[23][5] ), .QN(n903) );
  SDFFNSRXL \regfile_reg[23][4]  ( .D(n3030), .SI(n905), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4478), .Q(\regfile[23][4] ), .QN(n904) );
  SDFFNSRXL \regfile_reg[23][3]  ( .D(n3028), .SI(n906), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4478), .Q(\regfile[23][3] ), .QN(n905) );
  SDFFNSRXL \regfile_reg[23][2]  ( .D(n3026), .SI(n907), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4478), .Q(\regfile[23][2] ), .QN(n906) );
  SDFFNSRXL \regfile_reg[23][1]  ( .D(n3024), .SI(n908), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4478), .Q(\regfile[23][1] ), .QN(n907) );
  SDFFNSRXL \regfile_reg[23][0]  ( .D(n3022), .SI(n909), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4478), .Q(\regfile[23][0] ), .QN(n908) );
  SDFFNSRXL \regfile_reg[19][31]  ( .D(n2828), .SI(n1006), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4484), .Q(\regfile[19][31] ), .QN(n1005) );
  SDFFNSRXL \regfile_reg[19][30]  ( .D(n2826), .SI(n1007), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4484), .Q(\regfile[19][30] ), .QN(n1006) );
  SDFFNSRXL \regfile_reg[19][29]  ( .D(n2824), .SI(n1008), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4484), .Q(\regfile[19][29] ), .QN(n1007) );
  SDFFNSRXL \regfile_reg[19][28]  ( .D(n2822), .SI(n1009), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4484), .Q(\regfile[19][28] ), .QN(n1008) );
  SDFFNSRXL \regfile_reg[19][27]  ( .D(n2820), .SI(n1010), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4484), .Q(\regfile[19][27] ), .QN(n1009) );
  SDFFNSRXL \regfile_reg[19][26]  ( .D(n2818), .SI(n1011), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4484), .Q(\regfile[19][26] ), .QN(n1010) );
  SDFFNSRXL \regfile_reg[19][25]  ( .D(n2816), .SI(n1012), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4484), .Q(\regfile[19][25] ), .QN(n1011) );
  SDFFNSRXL \regfile_reg[19][24]  ( .D(n2814), .SI(n1013), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4484), .Q(\regfile[19][24] ), .QN(n1012) );
  SDFFNSRXL \regfile_reg[19][23]  ( .D(n2812), .SI(n1014), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4484), .Q(\regfile[19][23] ), .QN(n1013) );
  SDFFNSRXL \regfile_reg[19][22]  ( .D(n2810), .SI(n1015), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4484), .Q(\regfile[19][22] ), .QN(n1014) );
  SDFFNSRXL \regfile_reg[19][21]  ( .D(n2808), .SI(n1016), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4484), .Q(\regfile[19][21] ), .QN(n1015) );
  SDFFNSRXL \regfile_reg[19][20]  ( .D(n2806), .SI(n1017), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4484), .Q(\regfile[19][20] ), .QN(n1016) );
  SDFFNSRXL \regfile_reg[19][19]  ( .D(n2804), .SI(n1018), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4484), .Q(\regfile[19][19] ), .QN(n1017) );
  SDFFNSRXL \regfile_reg[19][18]  ( .D(n2802), .SI(n1019), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4484), .Q(\regfile[19][18] ), .QN(n1018) );
  SDFFNSRXL \regfile_reg[19][17]  ( .D(n2800), .SI(n1020), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4485), .Q(\regfile[19][17] ), .QN(n1019) );
  SDFFNSRXL \regfile_reg[19][16]  ( .D(n2798), .SI(n1021), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4485), .Q(\regfile[19][16] ), .QN(n1020) );
  SDFFNSRXL \regfile_reg[19][15]  ( .D(n2796), .SI(n1022), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4485), .Q(\regfile[19][15] ), .QN(n1021) );
  SDFFNSRXL \regfile_reg[19][14]  ( .D(n2794), .SI(n1023), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4485), .Q(\regfile[19][14] ), .QN(n1022) );
  SDFFNSRXL \regfile_reg[19][13]  ( .D(n2792), .SI(n1024), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4485), .Q(\regfile[19][13] ), .QN(n1023) );
  SDFFNSRXL \regfile_reg[19][12]  ( .D(n2790), .SI(n1025), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4485), .Q(\regfile[19][12] ), .QN(n1024) );
  SDFFNSRXL \regfile_reg[19][11]  ( .D(n2788), .SI(n1026), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4485), .Q(\regfile[19][11] ), .QN(n1025) );
  SDFFNSRXL \regfile_reg[19][10]  ( .D(n2786), .SI(n1027), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4485), .Q(\regfile[19][10] ), .QN(n1026) );
  SDFFNSRXL \regfile_reg[19][9]  ( .D(n2784), .SI(n1028), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4485), .Q(\regfile[19][9] ), .QN(n1027) );
  SDFFNSRXL \regfile_reg[19][8]  ( .D(n2782), .SI(n1029), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4485), .Q(\regfile[19][8] ), .QN(n1028) );
  SDFFNSRXL \regfile_reg[19][7]  ( .D(n2780), .SI(n1030), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4485), .Q(\regfile[19][7] ), .QN(n1029) );
  SDFFNSRXL \regfile_reg[19][6]  ( .D(n2778), .SI(n1031), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4485), .Q(\regfile[19][6] ), .QN(n1030) );
  SDFFNSRXL \regfile_reg[19][5]  ( .D(n2776), .SI(n1032), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4485), .Q(\regfile[19][5] ), .QN(n1031) );
  SDFFNSRXL \regfile_reg[19][4]  ( .D(n2774), .SI(n1033), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4485), .Q(\regfile[19][4] ), .QN(n1032) );
  SDFFNSRXL \regfile_reg[19][3]  ( .D(n2772), .SI(n1034), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4485), .Q(\regfile[19][3] ), .QN(n1033) );
  SDFFNSRXL \regfile_reg[19][2]  ( .D(n2770), .SI(n1035), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4485), .Q(\regfile[19][2] ), .QN(n1034) );
  SDFFNSRXL \regfile_reg[19][1]  ( .D(n2768), .SI(n1036), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4485), .Q(\regfile[19][1] ), .QN(n1035) );
  SDFFNSRXL \regfile_reg[19][0]  ( .D(n2766), .SI(n1037), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4485), .Q(\regfile[19][0] ), .QN(n1036) );
  SDFFNSRXL \regfile_reg[15][31]  ( .D(n2572), .SI(n1134), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4491), .Q(\regfile[15][31] ), .QN(n1133) );
  SDFFNSRXL \regfile_reg[15][30]  ( .D(n2570), .SI(n1135), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4491), .Q(\regfile[15][30] ), .QN(n1134) );
  SDFFNSRXL \regfile_reg[15][29]  ( .D(n2568), .SI(n1136), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4491), .Q(\regfile[15][29] ), .QN(n1135) );
  SDFFNSRXL \regfile_reg[15][28]  ( .D(n2566), .SI(n1137), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4491), .Q(\regfile[15][28] ), .QN(n1136) );
  SDFFNSRXL \regfile_reg[15][27]  ( .D(n2564), .SI(n1138), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4491), .Q(\regfile[15][27] ), .QN(n1137) );
  SDFFNSRXL \regfile_reg[15][26]  ( .D(n2562), .SI(n1139), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4491), .Q(\regfile[15][26] ), .QN(n1138) );
  SDFFNSRXL \regfile_reg[15][25]  ( .D(n2560), .SI(n1140), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4491), .Q(\regfile[15][25] ), .QN(n1139) );
  SDFFNSRXL \regfile_reg[15][24]  ( .D(n2558), .SI(n1141), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4491), .Q(\regfile[15][24] ), .QN(n1140) );
  SDFFNSRXL \regfile_reg[15][23]  ( .D(n2556), .SI(n1142), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4491), .Q(\regfile[15][23] ), .QN(n1141) );
  SDFFNSRXL \regfile_reg[15][22]  ( .D(n2554), .SI(n1143), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4491), .Q(\regfile[15][22] ), .QN(n1142) );
  SDFFNSRXL \regfile_reg[15][21]  ( .D(n2552), .SI(n1144), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4491), .Q(\regfile[15][21] ), .QN(n1143) );
  SDFFNSRXL \regfile_reg[15][20]  ( .D(n2550), .SI(n1145), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4491), .Q(\regfile[15][20] ), .QN(n1144) );
  SDFFNSRXL \regfile_reg[15][19]  ( .D(n2548), .SI(n1146), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4492), .Q(\regfile[15][19] ), .QN(n1145) );
  SDFFNSRXL \regfile_reg[15][18]  ( .D(n2546), .SI(n1147), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4492), .Q(\regfile[15][18] ), .QN(n1146) );
  SDFFNSRXL \regfile_reg[15][17]  ( .D(n2544), .SI(n1148), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4492), .Q(\regfile[15][17] ), .QN(n1147) );
  SDFFNSRXL \regfile_reg[15][16]  ( .D(n2542), .SI(n1149), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4492), .Q(\regfile[15][16] ), .QN(n1148) );
  SDFFNSRXL \regfile_reg[15][15]  ( .D(n2540), .SI(n1150), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4492), .Q(\regfile[15][15] ), .QN(n1149) );
  SDFFNSRXL \regfile_reg[15][14]  ( .D(n2538), .SI(n1151), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4492), .Q(\regfile[15][14] ), .QN(n1150) );
  SDFFNSRXL \regfile_reg[15][13]  ( .D(n2536), .SI(n1152), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4492), .Q(\regfile[15][13] ), .QN(n1151) );
  SDFFNSRXL \regfile_reg[15][12]  ( .D(n2534), .SI(n1153), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4492), .Q(\regfile[15][12] ), .QN(n1152) );
  SDFFNSRXL \regfile_reg[15][11]  ( .D(n2532), .SI(n1154), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4492), .Q(\regfile[15][11] ), .QN(n1153) );
  SDFFNSRXL \regfile_reg[15][10]  ( .D(n2530), .SI(n1155), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4492), .Q(\regfile[15][10] ), .QN(n1154) );
  SDFFNSRXL \regfile_reg[15][9]  ( .D(n2528), .SI(n1156), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4492), .Q(\regfile[15][9] ), .QN(n1155) );
  SDFFNSRXL \regfile_reg[15][8]  ( .D(n2526), .SI(n1157), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4492), .Q(\regfile[15][8] ), .QN(n1156) );
  SDFFNSRXL \regfile_reg[15][7]  ( .D(n2524), .SI(n1158), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4492), .Q(\regfile[15][7] ), .QN(n1157) );
  SDFFNSRXL \regfile_reg[15][6]  ( .D(n2522), .SI(n1159), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4492), .Q(\regfile[15][6] ), .QN(n1158) );
  SDFFNSRXL \regfile_reg[15][5]  ( .D(n2520), .SI(n1160), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4492), .Q(\regfile[15][5] ), .QN(n1159) );
  SDFFNSRXL \regfile_reg[15][4]  ( .D(n2518), .SI(n1161), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4492), .Q(\regfile[15][4] ), .QN(n1160) );
  SDFFNSRXL \regfile_reg[15][3]  ( .D(n2516), .SI(n1162), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4492), .Q(\regfile[15][3] ), .QN(n1161) );
  SDFFNSRXL \regfile_reg[15][2]  ( .D(n2514), .SI(n1163), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4492), .Q(\regfile[15][2] ), .QN(n1162) );
  SDFFNSRXL \regfile_reg[15][1]  ( .D(n2512), .SI(n1164), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4493), .Q(\regfile[15][1] ), .QN(n1163) );
  SDFFNSRXL \regfile_reg[15][0]  ( .D(n2510), .SI(n1165), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4493), .Q(\regfile[15][0] ), .QN(n1164) );
  SDFFNSRXL \regfile_reg[11][31]  ( .D(n2316), .SI(n1262), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4498), .Q(\regfile[11][31] ), .QN(n1261) );
  SDFFNSRXL \regfile_reg[11][30]  ( .D(n2314), .SI(n1263), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4498), .Q(\regfile[11][30] ), .QN(n1262) );
  SDFFNSRXL \regfile_reg[11][29]  ( .D(n2312), .SI(n1264), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4498), .Q(\regfile[11][29] ), .QN(n1263) );
  SDFFNSRXL \regfile_reg[11][28]  ( .D(n2310), .SI(n1265), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4498), .Q(\regfile[11][28] ), .QN(n1264) );
  SDFFNSRXL \regfile_reg[11][27]  ( .D(n2308), .SI(n1266), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4498), .Q(\regfile[11][27] ), .QN(n1265) );
  SDFFNSRXL \regfile_reg[11][26]  ( .D(n2306), .SI(n1267), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4498), .Q(\regfile[11][26] ), .QN(n1266) );
  SDFFNSRXL \regfile_reg[11][25]  ( .D(n2304), .SI(n1268), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4498), .Q(\regfile[11][25] ), .QN(n1267) );
  SDFFNSRXL \regfile_reg[11][24]  ( .D(n2302), .SI(n1269), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4498), .Q(\regfile[11][24] ), .QN(n1268) );
  SDFFNSRXL \regfile_reg[11][23]  ( .D(n2300), .SI(n1270), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4498), .Q(\regfile[11][23] ), .QN(n1269) );
  SDFFNSRXL \regfile_reg[11][22]  ( .D(n2298), .SI(n1271), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4498), .Q(\regfile[11][22] ), .QN(n1270) );
  SDFFNSRXL \regfile_reg[11][21]  ( .D(n2296), .SI(n1272), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4499), .Q(\regfile[11][21] ), .QN(n1271) );
  SDFFNSRXL \regfile_reg[11][20]  ( .D(n2294), .SI(n1273), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4499), .Q(\regfile[11][20] ), .QN(n1272) );
  SDFFNSRXL \regfile_reg[11][19]  ( .D(n2292), .SI(n1274), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4499), .Q(\regfile[11][19] ), .QN(n1273) );
  SDFFNSRXL \regfile_reg[11][18]  ( .D(n2290), .SI(n1275), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4499), .Q(\regfile[11][18] ), .QN(n1274) );
  SDFFNSRXL \regfile_reg[11][17]  ( .D(n2288), .SI(n1276), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4499), .Q(\regfile[11][17] ), .QN(n1275) );
  SDFFNSRXL \regfile_reg[11][16]  ( .D(n2286), .SI(n1277), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4499), .Q(\regfile[11][16] ), .QN(n1276) );
  SDFFNSRXL \regfile_reg[11][15]  ( .D(n2284), .SI(n1278), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4499), .Q(\regfile[11][15] ), .QN(n1277) );
  SDFFNSRXL \regfile_reg[11][14]  ( .D(n2282), .SI(n1279), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4499), .Q(\regfile[11][14] ), .QN(n1278) );
  SDFFNSRXL \regfile_reg[11][13]  ( .D(n2280), .SI(n1280), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4499), .Q(\regfile[11][13] ), .QN(n1279) );
  SDFFNSRXL \regfile_reg[11][12]  ( .D(n2278), .SI(n1281), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4499), .Q(\regfile[11][12] ), .QN(n1280) );
  SDFFNSRXL \regfile_reg[11][11]  ( .D(n2276), .SI(n1282), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4499), .Q(\regfile[11][11] ), .QN(n1281) );
  SDFFNSRXL \regfile_reg[11][10]  ( .D(n2274), .SI(n1283), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4499), .Q(\regfile[11][10] ), .QN(n1282) );
  SDFFNSRXL \regfile_reg[11][9]  ( .D(n2272), .SI(n1284), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4499), .Q(\regfile[11][9] ), .QN(n1283) );
  SDFFNSRXL \regfile_reg[11][8]  ( .D(n2270), .SI(n1285), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4499), .Q(\regfile[11][8] ), .QN(n1284) );
  SDFFNSRXL \regfile_reg[11][7]  ( .D(n2268), .SI(n1286), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4499), .Q(\regfile[11][7] ), .QN(n1285) );
  SDFFNSRXL \regfile_reg[11][6]  ( .D(n2266), .SI(n1287), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4499), .Q(\regfile[11][6] ), .QN(n1286) );
  SDFFNSRXL \regfile_reg[11][5]  ( .D(n2264), .SI(n1288), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4499), .Q(\regfile[11][5] ), .QN(n1287) );
  SDFFNSRXL \regfile_reg[11][4]  ( .D(n2262), .SI(n1289), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4499), .Q(\regfile[11][4] ), .QN(n1288) );
  SDFFNSRXL \regfile_reg[11][3]  ( .D(n2260), .SI(n1290), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4500), .Q(\regfile[11][3] ), .QN(n1289) );
  SDFFNSRXL \regfile_reg[11][2]  ( .D(n2258), .SI(n1291), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4500), .Q(\regfile[11][2] ), .QN(n1290) );
  SDFFNSRXL \regfile_reg[11][1]  ( .D(n2256), .SI(n1292), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4500), .Q(\regfile[11][1] ), .QN(n1291) );
  SDFFNSRXL \regfile_reg[11][0]  ( .D(n2254), .SI(n1293), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4500), .Q(\regfile[11][0] ), .QN(n1292) );
  SDFFNSRXL \regfile_reg[7][31]  ( .D(n2060), .SI(n1390), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4505), .Q(\regfile[7][31] ), .QN(n1389) );
  SDFFNSRXL \regfile_reg[7][30]  ( .D(n2058), .SI(n1391), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4505), .Q(\regfile[7][30] ), .QN(n1390) );
  SDFFNSRXL \regfile_reg[7][29]  ( .D(n2056), .SI(n1392), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4505), .Q(\regfile[7][29] ), .QN(n1391) );
  SDFFNSRXL \regfile_reg[7][28]  ( .D(n2054), .SI(n1393), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4505), .Q(\regfile[7][28] ), .QN(n1392) );
  SDFFNSRXL \regfile_reg[7][27]  ( .D(n2052), .SI(n1394), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4505), .Q(\regfile[7][27] ), .QN(n1393) );
  SDFFNSRXL \regfile_reg[7][26]  ( .D(n2050), .SI(n1395), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4505), .Q(\regfile[7][26] ), .QN(n1394) );
  SDFFNSRXL \regfile_reg[7][25]  ( .D(n2048), .SI(n1396), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4505), .Q(\regfile[7][25] ), .QN(n1395) );
  SDFFNSRXL \regfile_reg[7][24]  ( .D(n2046), .SI(n1397), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4505), .Q(\regfile[7][24] ), .QN(n1396) );
  SDFFNSRXL \regfile_reg[7][23]  ( .D(n2044), .SI(n1398), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4506), .Q(\regfile[7][23] ), .QN(n1397) );
  SDFFNSRXL \regfile_reg[7][22]  ( .D(n2042), .SI(n1399), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4506), .Q(\regfile[7][22] ), .QN(n1398) );
  SDFFNSRXL \regfile_reg[7][21]  ( .D(n2040), .SI(n1400), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4506), .Q(\regfile[7][21] ), .QN(n1399) );
  SDFFNSRXL \regfile_reg[7][20]  ( .D(n2038), .SI(n1401), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4506), .Q(\regfile[7][20] ), .QN(n1400) );
  SDFFNSRXL \regfile_reg[7][19]  ( .D(n2036), .SI(n1402), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4506), .Q(\regfile[7][19] ), .QN(n1401) );
  SDFFNSRXL \regfile_reg[7][18]  ( .D(n2034), .SI(n1403), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4506), .Q(\regfile[7][18] ), .QN(n1402) );
  SDFFNSRXL \regfile_reg[7][17]  ( .D(n2032), .SI(n1404), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4506), .Q(\regfile[7][17] ), .QN(n1403) );
  SDFFNSRXL \regfile_reg[7][16]  ( .D(n2030), .SI(n1405), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4506), .Q(\regfile[7][16] ), .QN(n1404) );
  SDFFNSRXL \regfile_reg[7][15]  ( .D(n2028), .SI(n1406), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4506), .Q(\regfile[7][15] ), .QN(n1405) );
  SDFFNSRXL \regfile_reg[7][14]  ( .D(n2026), .SI(n1407), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4506), .Q(\regfile[7][14] ), .QN(n1406) );
  SDFFNSRXL \regfile_reg[7][13]  ( .D(n2024), .SI(n1408), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4506), .Q(\regfile[7][13] ), .QN(n1407) );
  SDFFNSRXL \regfile_reg[7][12]  ( .D(n2022), .SI(n1409), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4506), .Q(\regfile[7][12] ), .QN(n1408) );
  SDFFNSRXL \regfile_reg[7][11]  ( .D(n2020), .SI(n1410), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4506), .Q(\regfile[7][11] ), .QN(n1409) );
  SDFFNSRXL \regfile_reg[7][10]  ( .D(n2018), .SI(n1411), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4506), .Q(\regfile[7][10] ), .QN(n1410) );
  SDFFNSRXL \regfile_reg[7][9]  ( .D(n2016), .SI(n1412), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4506), .Q(\regfile[7][9] ), .QN(n1411) );
  SDFFNSRXL \regfile_reg[7][8]  ( .D(n2014), .SI(n1413), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4506), .Q(\regfile[7][8] ), .QN(n1412) );
  SDFFNSRXL \regfile_reg[7][7]  ( .D(n2012), .SI(n1414), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4506), .Q(\regfile[7][7] ), .QN(n1413) );
  SDFFNSRXL \regfile_reg[7][6]  ( .D(n2010), .SI(n1415), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4506), .Q(\regfile[7][6] ), .QN(n1414) );
  SDFFNSRXL \regfile_reg[7][5]  ( .D(n2008), .SI(n1416), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4507), .Q(\regfile[7][5] ), .QN(n1415) );
  SDFFNSRXL \regfile_reg[7][4]  ( .D(n2006), .SI(n1417), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4507), .Q(\regfile[7][4] ), .QN(n1416) );
  SDFFNSRXL \regfile_reg[7][3]  ( .D(n2004), .SI(n1418), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4507), .Q(\regfile[7][3] ), .QN(n1417) );
  SDFFNSRXL \regfile_reg[7][2]  ( .D(n2002), .SI(n1419), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4507), .Q(\regfile[7][2] ), .QN(n1418) );
  SDFFNSRXL \regfile_reg[7][1]  ( .D(n2000), .SI(n1420), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4507), .Q(\regfile[7][1] ), .QN(n1419) );
  SDFFNSRXL \regfile_reg[7][0]  ( .D(n1998), .SI(n1421), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4507), .Q(\regfile[7][0] ), .QN(n1420) );
  SDFFNSRXL \regfile_reg[29][31]  ( .D(n3468), .SI(n686), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4466), .Q(\regfile[29][31] ), .QN(n685) );
  SDFFNSRXL \regfile_reg[29][30]  ( .D(n3466), .SI(n687), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4466), .Q(\regfile[29][30] ), .QN(n686) );
  SDFFNSRXL \regfile_reg[29][29]  ( .D(n3464), .SI(n688), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4466), .Q(\regfile[29][29] ), .QN(n687) );
  SDFFNSRXL \regfile_reg[29][28]  ( .D(n3462), .SI(n689), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4466), .Q(\regfile[29][28] ), .QN(n688) );
  SDFFNSRXL \regfile_reg[29][27]  ( .D(n3460), .SI(n690), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4466), .Q(\regfile[29][27] ), .QN(n689) );
  SDFFNSRXL \regfile_reg[29][26]  ( .D(n3458), .SI(n691), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4466), .Q(\regfile[29][26] ), .QN(n690) );
  SDFFNSRXL \regfile_reg[29][25]  ( .D(n3456), .SI(n692), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4466), .Q(\regfile[29][25] ), .QN(n691) );
  SDFFNSRXL \regfile_reg[29][24]  ( .D(n3454), .SI(n693), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4466), .Q(\regfile[29][24] ), .QN(n692) );
  SDFFNSRXL \regfile_reg[29][23]  ( .D(n3452), .SI(n694), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4466), .Q(\regfile[29][23] ), .QN(n693) );
  SDFFNSRXL \regfile_reg[29][22]  ( .D(n3450), .SI(n695), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4466), .Q(\regfile[29][22] ), .QN(n694) );
  SDFFNSRXL \regfile_reg[29][21]  ( .D(n3448), .SI(n696), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4467), .Q(\regfile[29][21] ), .QN(n695) );
  SDFFNSRXL \regfile_reg[29][20]  ( .D(n3446), .SI(n697), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4467), .Q(\regfile[29][20] ), .QN(n696) );
  SDFFNSRXL \regfile_reg[29][19]  ( .D(n3444), .SI(n698), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4467), .Q(\regfile[29][19] ), .QN(n697) );
  SDFFNSRXL \regfile_reg[29][18]  ( .D(n3442), .SI(n699), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4467), .Q(\regfile[29][18] ), .QN(n698) );
  SDFFNSRXL \regfile_reg[29][17]  ( .D(n3440), .SI(n700), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4467), .Q(\regfile[29][17] ), .QN(n699) );
  SDFFNSRXL \regfile_reg[29][16]  ( .D(n3438), .SI(n701), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4467), .Q(\regfile[29][16] ), .QN(n700) );
  SDFFNSRXL \regfile_reg[29][15]  ( .D(n3436), .SI(n702), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4467), .Q(\regfile[29][15] ), .QN(n701) );
  SDFFNSRXL \regfile_reg[29][14]  ( .D(n3434), .SI(n703), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4467), .Q(\regfile[29][14] ), .QN(n702) );
  SDFFNSRXL \regfile_reg[29][13]  ( .D(n3432), .SI(n704), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4467), .Q(\regfile[29][13] ), .QN(n703) );
  SDFFNSRXL \regfile_reg[29][12]  ( .D(n3430), .SI(n705), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4467), .Q(\regfile[29][12] ), .QN(n704) );
  SDFFNSRXL \regfile_reg[29][11]  ( .D(n3428), .SI(n706), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4467), .Q(\regfile[29][11] ), .QN(n705) );
  SDFFNSRXL \regfile_reg[29][10]  ( .D(n3426), .SI(n707), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4467), .Q(\regfile[29][10] ), .QN(n706) );
  SDFFNSRXL \regfile_reg[29][9]  ( .D(n3424), .SI(n708), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4467), .Q(\regfile[29][9] ), .QN(n707) );
  SDFFNSRXL \regfile_reg[29][8]  ( .D(n3422), .SI(n709), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4467), .Q(\regfile[29][8] ), .QN(n708) );
  SDFFNSRXL \regfile_reg[29][7]  ( .D(n3420), .SI(n710), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4467), .Q(\regfile[29][7] ), .QN(n709) );
  SDFFNSRXL \regfile_reg[29][6]  ( .D(n3418), .SI(n711), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4467), .Q(\regfile[29][6] ), .QN(n710) );
  SDFFNSRXL \regfile_reg[29][5]  ( .D(n3416), .SI(n712), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4467), .Q(\regfile[29][5] ), .QN(n711) );
  SDFFNSRXL \regfile_reg[29][4]  ( .D(n3414), .SI(n713), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4467), .Q(\regfile[29][4] ), .QN(n712) );
  SDFFNSRXL \regfile_reg[29][3]  ( .D(n3412), .SI(n714), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4468), .Q(\regfile[29][3] ), .QN(n713) );
  SDFFNSRXL \regfile_reg[29][2]  ( .D(n3410), .SI(n715), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4468), .Q(\regfile[29][2] ), .QN(n714) );
  SDFFNSRXL \regfile_reg[29][1]  ( .D(n3408), .SI(n716), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4468), .Q(\regfile[29][1] ), .QN(n715) );
  SDFFNSRXL \regfile_reg[29][0]  ( .D(n3406), .SI(n717), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4468), .Q(\regfile[29][0] ), .QN(n716) );
  SDFFNSRXL \regfile_reg[25][31]  ( .D(n3212), .SI(n814), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4473), .Q(\regfile[25][31] ), .QN(n813) );
  SDFFNSRXL \regfile_reg[25][30]  ( .D(n3210), .SI(n815), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4473), .Q(\regfile[25][30] ), .QN(n814) );
  SDFFNSRXL \regfile_reg[25][29]  ( .D(n3208), .SI(n816), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4473), .Q(\regfile[25][29] ), .QN(n815) );
  SDFFNSRXL \regfile_reg[25][28]  ( .D(n3206), .SI(n817), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4473), .Q(\regfile[25][28] ), .QN(n816) );
  SDFFNSRXL \regfile_reg[25][27]  ( .D(n3204), .SI(n818), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4473), .Q(\regfile[25][27] ), .QN(n817) );
  SDFFNSRXL \regfile_reg[25][26]  ( .D(n3202), .SI(n819), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4473), .Q(\regfile[25][26] ), .QN(n818) );
  SDFFNSRXL \regfile_reg[25][25]  ( .D(n3200), .SI(n820), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4473), .Q(\regfile[25][25] ), .QN(n819) );
  SDFFNSRXL \regfile_reg[25][24]  ( .D(n3198), .SI(n821), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4473), .Q(\regfile[25][24] ), .QN(n820) );
  SDFFNSRXL \regfile_reg[25][23]  ( .D(n3196), .SI(n822), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4474), .Q(\regfile[25][23] ), .QN(n821) );
  SDFFNSRXL \regfile_reg[25][22]  ( .D(n3194), .SI(n823), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4474), .Q(\regfile[25][22] ), .QN(n822) );
  SDFFNSRXL \regfile_reg[25][21]  ( .D(n3192), .SI(n824), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4474), .Q(\regfile[25][21] ), .QN(n823) );
  SDFFNSRXL \regfile_reg[25][20]  ( .D(n3190), .SI(n825), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4474), .Q(\regfile[25][20] ), .QN(n824) );
  SDFFNSRXL \regfile_reg[25][19]  ( .D(n3188), .SI(n826), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4474), .Q(\regfile[25][19] ), .QN(n825) );
  SDFFNSRXL \regfile_reg[25][18]  ( .D(n3186), .SI(n827), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4474), .Q(\regfile[25][18] ), .QN(n826) );
  SDFFNSRXL \regfile_reg[25][17]  ( .D(n3184), .SI(n828), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4474), .Q(\regfile[25][17] ), .QN(n827) );
  SDFFNSRXL \regfile_reg[25][16]  ( .D(n3182), .SI(n829), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4474), .Q(\regfile[25][16] ), .QN(n828) );
  SDFFNSRXL \regfile_reg[25][15]  ( .D(n3180), .SI(n830), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4474), .Q(\regfile[25][15] ), .QN(n829) );
  SDFFNSRXL \regfile_reg[25][14]  ( .D(n3178), .SI(n831), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4474), .Q(\regfile[25][14] ), .QN(n830) );
  SDFFNSRXL \regfile_reg[25][13]  ( .D(n3176), .SI(n832), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4474), .Q(\regfile[25][13] ), .QN(n831) );
  SDFFNSRXL \regfile_reg[25][12]  ( .D(n3174), .SI(n833), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4474), .Q(\regfile[25][12] ), .QN(n832) );
  SDFFNSRXL \regfile_reg[25][11]  ( .D(n3172), .SI(n834), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4474), .Q(\regfile[25][11] ), .QN(n833) );
  SDFFNSRXL \regfile_reg[25][10]  ( .D(n3170), .SI(n835), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4474), .Q(\regfile[25][10] ), .QN(n834) );
  SDFFNSRXL \regfile_reg[25][9]  ( .D(n3168), .SI(n836), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4474), .Q(\regfile[25][9] ), .QN(n835) );
  SDFFNSRXL \regfile_reg[25][8]  ( .D(n3166), .SI(n837), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4474), .Q(\regfile[25][8] ), .QN(n836) );
  SDFFNSRXL \regfile_reg[25][7]  ( .D(n3164), .SI(n838), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4474), .Q(\regfile[25][7] ), .QN(n837) );
  SDFFNSRXL \regfile_reg[25][6]  ( .D(n3162), .SI(n839), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4474), .Q(\regfile[25][6] ), .QN(n838) );
  SDFFNSRXL \regfile_reg[25][5]  ( .D(n3160), .SI(n840), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4475), .Q(\regfile[25][5] ), .QN(n839) );
  SDFFNSRXL \regfile_reg[25][4]  ( .D(n3158), .SI(n841), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4475), .Q(\regfile[25][4] ), .QN(n840) );
  SDFFNSRXL \regfile_reg[25][3]  ( .D(n3156), .SI(n842), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4475), .Q(\regfile[25][3] ), .QN(n841) );
  SDFFNSRXL \regfile_reg[25][2]  ( .D(n3154), .SI(n843), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4475), .Q(\regfile[25][2] ), .QN(n842) );
  SDFFNSRXL \regfile_reg[25][1]  ( .D(n3152), .SI(n844), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4475), .Q(\regfile[25][1] ), .QN(n843) );
  SDFFNSRXL \regfile_reg[25][0]  ( .D(n3150), .SI(n845), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4475), .Q(\regfile[25][0] ), .QN(n844) );
  SDFFNSRXL \regfile_reg[21][31]  ( .D(n2956), .SI(n942), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4480), .Q(\regfile[21][31] ), .QN(n941) );
  SDFFNSRXL \regfile_reg[21][30]  ( .D(n2954), .SI(n943), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4480), .Q(\regfile[21][30] ), .QN(n942) );
  SDFFNSRXL \regfile_reg[21][29]  ( .D(n2952), .SI(n944), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4480), .Q(\regfile[21][29] ), .QN(n943) );
  SDFFNSRXL \regfile_reg[21][28]  ( .D(n2950), .SI(n945), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4480), .Q(\regfile[21][28] ), .QN(n944) );
  SDFFNSRXL \regfile_reg[21][27]  ( .D(n2948), .SI(n946), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4480), .Q(\regfile[21][27] ), .QN(n945) );
  SDFFNSRXL \regfile_reg[21][26]  ( .D(n2946), .SI(n947), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4480), .Q(\regfile[21][26] ), .QN(n946) );
  SDFFNSRXL \regfile_reg[21][25]  ( .D(n2944), .SI(n948), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4481), .Q(\regfile[21][25] ), .QN(n947) );
  SDFFNSRXL \regfile_reg[21][24]  ( .D(n2942), .SI(n949), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4481), .Q(\regfile[21][24] ), .QN(n948) );
  SDFFNSRXL \regfile_reg[21][23]  ( .D(n2940), .SI(n950), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4481), .Q(\regfile[21][23] ), .QN(n949) );
  SDFFNSRXL \regfile_reg[21][22]  ( .D(n2938), .SI(n951), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4481), .Q(\regfile[21][22] ), .QN(n950) );
  SDFFNSRXL \regfile_reg[21][21]  ( .D(n2936), .SI(n952), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4481), .Q(\regfile[21][21] ), .QN(n951) );
  SDFFNSRXL \regfile_reg[21][20]  ( .D(n2934), .SI(n953), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4481), .Q(\regfile[21][20] ), .QN(n952) );
  SDFFNSRXL \regfile_reg[21][19]  ( .D(n2932), .SI(n954), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4481), .Q(\regfile[21][19] ), .QN(n953) );
  SDFFNSRXL \regfile_reg[21][18]  ( .D(n2930), .SI(n955), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4481), .Q(\regfile[21][18] ), .QN(n954) );
  SDFFNSRXL \regfile_reg[21][17]  ( .D(n2928), .SI(n956), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4481), .Q(\regfile[21][17] ), .QN(n955) );
  SDFFNSRXL \regfile_reg[21][16]  ( .D(n2926), .SI(n957), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4481), .Q(\regfile[21][16] ), .QN(n956) );
  SDFFNSRXL \regfile_reg[21][15]  ( .D(n2924), .SI(n958), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4481), .Q(\regfile[21][15] ), .QN(n957) );
  SDFFNSRXL \regfile_reg[21][14]  ( .D(n2922), .SI(n959), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4481), .Q(\regfile[21][14] ), .QN(n958) );
  SDFFNSRXL \regfile_reg[21][13]  ( .D(n2920), .SI(n960), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4481), .Q(\regfile[21][13] ), .QN(n959) );
  SDFFNSRXL \regfile_reg[21][12]  ( .D(n2918), .SI(n961), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4481), .Q(\regfile[21][12] ), .QN(n960) );
  SDFFNSRXL \regfile_reg[21][11]  ( .D(n2916), .SI(n962), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4481), .Q(\regfile[21][11] ), .QN(n961) );
  SDFFNSRXL \regfile_reg[21][10]  ( .D(n2914), .SI(n963), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4481), .Q(\regfile[21][10] ), .QN(n962) );
  SDFFNSRXL \regfile_reg[21][9]  ( .D(n2912), .SI(n964), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4481), .Q(\regfile[21][9] ), .QN(n963) );
  SDFFNSRXL \regfile_reg[21][8]  ( .D(n2910), .SI(n965), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4481), .Q(\regfile[21][8] ), .QN(n964) );
  SDFFNSRXL \regfile_reg[21][7]  ( .D(n2908), .SI(n966), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4482), .Q(\regfile[21][7] ), .QN(n965) );
  SDFFNSRXL \regfile_reg[21][6]  ( .D(n2906), .SI(n967), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4482), .Q(\regfile[21][6] ), .QN(n966) );
  SDFFNSRXL \regfile_reg[21][5]  ( .D(n2904), .SI(n968), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4482), .Q(\regfile[21][5] ), .QN(n967) );
  SDFFNSRXL \regfile_reg[21][4]  ( .D(n2902), .SI(n969), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4482), .Q(\regfile[21][4] ), .QN(n968) );
  SDFFNSRXL \regfile_reg[21][3]  ( .D(n2900), .SI(n970), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4482), .Q(\regfile[21][3] ), .QN(n969) );
  SDFFNSRXL \regfile_reg[21][2]  ( .D(n2898), .SI(n971), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4482), .Q(\regfile[21][2] ), .QN(n970) );
  SDFFNSRXL \regfile_reg[21][1]  ( .D(n2896), .SI(n972), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4482), .Q(\regfile[21][1] ), .QN(n971) );
  SDFFNSRXL \regfile_reg[21][0]  ( .D(n2894), .SI(n973), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4482), .Q(\regfile[21][0] ), .QN(n972) );
  SDFFNSRXL \regfile_reg[17][31]  ( .D(n2700), .SI(n1070), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4487), .Q(\regfile[17][31] ), .QN(n1069) );
  SDFFNSRXL \regfile_reg[17][30]  ( .D(n2698), .SI(n1071), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4487), .Q(\regfile[17][30] ), .QN(n1070) );
  SDFFNSRXL \regfile_reg[17][29]  ( .D(n2696), .SI(n1072), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4487), .Q(\regfile[17][29] ), .QN(n1071) );
  SDFFNSRXL \regfile_reg[17][28]  ( .D(n2694), .SI(n1073), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4487), .Q(\regfile[17][28] ), .QN(n1072) );
  SDFFNSRXL \regfile_reg[17][27]  ( .D(n2692), .SI(n1074), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4488), .Q(\regfile[17][27] ), .QN(n1073) );
  SDFFNSRXL \regfile_reg[17][26]  ( .D(n2690), .SI(n1075), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4488), .Q(\regfile[17][26] ), .QN(n1074) );
  SDFFNSRXL \regfile_reg[17][25]  ( .D(n2688), .SI(n1076), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4488), .Q(\regfile[17][25] ), .QN(n1075) );
  SDFFNSRXL \regfile_reg[17][24]  ( .D(n2686), .SI(n1077), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4488), .Q(\regfile[17][24] ), .QN(n1076) );
  SDFFNSRXL \regfile_reg[17][23]  ( .D(n2684), .SI(n1078), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4488), .Q(\regfile[17][23] ), .QN(n1077) );
  SDFFNSRXL \regfile_reg[17][22]  ( .D(n2682), .SI(n1079), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4488), .Q(\regfile[17][22] ), .QN(n1078) );
  SDFFNSRXL \regfile_reg[17][21]  ( .D(n2680), .SI(n1080), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4488), .Q(\regfile[17][21] ), .QN(n1079) );
  SDFFNSRXL \regfile_reg[17][20]  ( .D(n2678), .SI(n1081), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4488), .Q(\regfile[17][20] ), .QN(n1080) );
  SDFFNSRXL \regfile_reg[17][19]  ( .D(n2676), .SI(n1082), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4488), .Q(\regfile[17][19] ), .QN(n1081) );
  SDFFNSRXL \regfile_reg[17][18]  ( .D(n2674), .SI(n1083), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4488), .Q(\regfile[17][18] ), .QN(n1082) );
  SDFFNSRXL \regfile_reg[17][17]  ( .D(n2672), .SI(n1084), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4488), .Q(\regfile[17][17] ), .QN(n1083) );
  SDFFNSRXL \regfile_reg[17][16]  ( .D(n2670), .SI(n1085), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4488), .Q(\regfile[17][16] ), .QN(n1084) );
  SDFFNSRXL \regfile_reg[17][15]  ( .D(n2668), .SI(n1086), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4488), .Q(\regfile[17][15] ), .QN(n1085) );
  SDFFNSRXL \regfile_reg[17][14]  ( .D(n2666), .SI(n1087), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4488), .Q(\regfile[17][14] ), .QN(n1086) );
  SDFFNSRXL \regfile_reg[17][13]  ( .D(n2664), .SI(n1088), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4488), .Q(\regfile[17][13] ), .QN(n1087) );
  SDFFNSRXL \regfile_reg[17][12]  ( .D(n2662), .SI(n1089), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4488), .Q(\regfile[17][12] ), .QN(n1088) );
  SDFFNSRXL \regfile_reg[17][11]  ( .D(n2660), .SI(n1090), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4488), .Q(\regfile[17][11] ), .QN(n1089) );
  SDFFNSRXL \regfile_reg[17][10]  ( .D(n2658), .SI(n1091), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4488), .Q(\regfile[17][10] ), .QN(n1090) );
  SDFFNSRXL \regfile_reg[17][9]  ( .D(n2656), .SI(n1092), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4489), .Q(\regfile[17][9] ), .QN(n1091) );
  SDFFNSRXL \regfile_reg[17][8]  ( .D(n2654), .SI(n1093), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4489), .Q(\regfile[17][8] ), .QN(n1092) );
  SDFFNSRXL \regfile_reg[17][7]  ( .D(n2652), .SI(n1094), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4489), .Q(\regfile[17][7] ), .QN(n1093) );
  SDFFNSRXL \regfile_reg[17][6]  ( .D(n2650), .SI(n1095), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4489), .Q(\regfile[17][6] ), .QN(n1094) );
  SDFFNSRXL \regfile_reg[17][5]  ( .D(n2648), .SI(n1096), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4489), .Q(\regfile[17][5] ), .QN(n1095) );
  SDFFNSRXL \regfile_reg[17][4]  ( .D(n2646), .SI(n1097), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4489), .Q(\regfile[17][4] ), .QN(n1096) );
  SDFFNSRXL \regfile_reg[17][3]  ( .D(n2644), .SI(n1098), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4489), .Q(\regfile[17][3] ), .QN(n1097) );
  SDFFNSRXL \regfile_reg[17][2]  ( .D(n2642), .SI(n1099), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4489), .Q(\regfile[17][2] ), .QN(n1098) );
  SDFFNSRXL \regfile_reg[17][1]  ( .D(n2640), .SI(n1100), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4489), .Q(\regfile[17][1] ), .QN(n1099) );
  SDFFNSRXL \regfile_reg[17][0]  ( .D(n2638), .SI(n1101), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4489), .Q(\regfile[17][0] ), .QN(n1100) );
  SDFFNSRXL \regfile_reg[13][31]  ( .D(n2444), .SI(n1198), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4494), .Q(\regfile[13][31] ), .QN(n1197) );
  SDFFNSRXL \regfile_reg[13][30]  ( .D(n2442), .SI(n1199), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4494), .Q(\regfile[13][30] ), .QN(n1198) );
  SDFFNSRXL \regfile_reg[13][29]  ( .D(n2440), .SI(n1200), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4495), .Q(\regfile[13][29] ), .QN(n1199) );
  SDFFNSRXL \regfile_reg[13][28]  ( .D(n2438), .SI(n1201), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4495), .Q(\regfile[13][28] ), .QN(n1200) );
  SDFFNSRXL \regfile_reg[13][27]  ( .D(n2436), .SI(n1202), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4495), .Q(\regfile[13][27] ), .QN(n1201) );
  SDFFNSRXL \regfile_reg[13][26]  ( .D(n2434), .SI(n1203), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4495), .Q(\regfile[13][26] ), .QN(n1202) );
  SDFFNSRXL \regfile_reg[13][25]  ( .D(n2432), .SI(n1204), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4495), .Q(\regfile[13][25] ), .QN(n1203) );
  SDFFNSRXL \regfile_reg[13][24]  ( .D(n2430), .SI(n1205), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4495), .Q(\regfile[13][24] ), .QN(n1204) );
  SDFFNSRXL \regfile_reg[13][23]  ( .D(n2428), .SI(n1206), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4495), .Q(\regfile[13][23] ), .QN(n1205) );
  SDFFNSRXL \regfile_reg[13][22]  ( .D(n2426), .SI(n1207), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4495), .Q(\regfile[13][22] ), .QN(n1206) );
  SDFFNSRXL \regfile_reg[13][21]  ( .D(n2424), .SI(n1208), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4495), .Q(\regfile[13][21] ), .QN(n1207) );
  SDFFNSRXL \regfile_reg[13][20]  ( .D(n2422), .SI(n1209), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4495), .Q(\regfile[13][20] ), .QN(n1208) );
  SDFFNSRXL \regfile_reg[13][19]  ( .D(n2420), .SI(n1210), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4495), .Q(\regfile[13][19] ), .QN(n1209) );
  SDFFNSRXL \regfile_reg[13][18]  ( .D(n2418), .SI(n1211), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4495), .Q(\regfile[13][18] ), .QN(n1210) );
  SDFFNSRXL \regfile_reg[13][17]  ( .D(n2416), .SI(n1212), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4495), .Q(\regfile[13][17] ), .QN(n1211) );
  SDFFNSRXL \regfile_reg[13][16]  ( .D(n2414), .SI(n1213), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4495), .Q(\regfile[13][16] ), .QN(n1212) );
  SDFFNSRXL \regfile_reg[13][15]  ( .D(n2412), .SI(n1214), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4495), .Q(\regfile[13][15] ), .QN(n1213) );
  SDFFNSRXL \regfile_reg[13][14]  ( .D(n2410), .SI(n1215), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4495), .Q(\regfile[13][14] ), .QN(n1214) );
  SDFFNSRXL \regfile_reg[13][13]  ( .D(n2408), .SI(n1216), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4495), .Q(\regfile[13][13] ), .QN(n1215) );
  SDFFNSRXL \regfile_reg[13][12]  ( .D(n2406), .SI(n1217), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4495), .Q(\regfile[13][12] ), .QN(n1216) );
  SDFFNSRXL \regfile_reg[13][11]  ( .D(n2404), .SI(n1218), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4496), .Q(\regfile[13][11] ), .QN(n1217) );
  SDFFNSRXL \regfile_reg[13][10]  ( .D(n2402), .SI(n1219), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4496), .Q(\regfile[13][10] ), .QN(n1218) );
  SDFFNSRXL \regfile_reg[13][9]  ( .D(n2400), .SI(n1220), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4496), .Q(\regfile[13][9] ), .QN(n1219) );
  SDFFNSRXL \regfile_reg[13][8]  ( .D(n2398), .SI(n1221), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4496), .Q(\regfile[13][8] ), .QN(n1220) );
  SDFFNSRXL \regfile_reg[13][7]  ( .D(n2396), .SI(n1222), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4496), .Q(\regfile[13][7] ), .QN(n1221) );
  SDFFNSRXL \regfile_reg[13][6]  ( .D(n2394), .SI(n1223), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4496), .Q(\regfile[13][6] ), .QN(n1222) );
  SDFFNSRXL \regfile_reg[13][5]  ( .D(n2392), .SI(n1224), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4496), .Q(\regfile[13][5] ), .QN(n1223) );
  SDFFNSRXL \regfile_reg[13][4]  ( .D(n2390), .SI(n1225), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4496), .Q(\regfile[13][4] ), .QN(n1224) );
  SDFFNSRXL \regfile_reg[13][3]  ( .D(n2388), .SI(n1226), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4496), .Q(\regfile[13][3] ), .QN(n1225) );
  SDFFNSRXL \regfile_reg[13][2]  ( .D(n2386), .SI(n1227), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4496), .Q(\regfile[13][2] ), .QN(n1226) );
  SDFFNSRXL \regfile_reg[13][1]  ( .D(n2384), .SI(n1228), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4496), .Q(\regfile[13][1] ), .QN(n1227) );
  SDFFNSRXL \regfile_reg[13][0]  ( .D(n2382), .SI(n1229), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4496), .Q(\regfile[13][0] ), .QN(n1228) );
  SDFFNSRXL \regfile_reg[9][31]  ( .D(n2188), .SI(n1326), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4502), .Q(\regfile[9][31] ), .QN(n1325) );
  SDFFNSRXL \regfile_reg[9][30]  ( .D(n2186), .SI(n1327), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4502), .Q(\regfile[9][30] ), .QN(n1326) );
  SDFFNSRXL \regfile_reg[9][29]  ( .D(n2184), .SI(n1328), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4502), .Q(\regfile[9][29] ), .QN(n1327) );
  SDFFNSRXL \regfile_reg[9][28]  ( .D(n2182), .SI(n1329), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4502), .Q(\regfile[9][28] ), .QN(n1328) );
  SDFFNSRXL \regfile_reg[9][27]  ( .D(n2180), .SI(n1330), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4502), .Q(\regfile[9][27] ), .QN(n1329) );
  SDFFNSRXL \regfile_reg[9][26]  ( .D(n2178), .SI(n1331), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4502), .Q(\regfile[9][26] ), .QN(n1330) );
  SDFFNSRXL \regfile_reg[9][25]  ( .D(n2176), .SI(n1332), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4502), .Q(\regfile[9][25] ), .QN(n1331) );
  SDFFNSRXL \regfile_reg[9][24]  ( .D(n2174), .SI(n1333), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4502), .Q(\regfile[9][24] ), .QN(n1332) );
  SDFFNSRXL \regfile_reg[9][23]  ( .D(n2172), .SI(n1334), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4502), .Q(\regfile[9][23] ), .QN(n1333) );
  SDFFNSRXL \regfile_reg[9][22]  ( .D(n2170), .SI(n1335), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4502), .Q(\regfile[9][22] ), .QN(n1334) );
  SDFFNSRXL \regfile_reg[9][21]  ( .D(n2168), .SI(n1336), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4502), .Q(\regfile[9][21] ), .QN(n1335) );
  SDFFNSRXL \regfile_reg[9][20]  ( .D(n2166), .SI(n1337), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4502), .Q(\regfile[9][20] ), .QN(n1336) );
  SDFFNSRXL \regfile_reg[9][19]  ( .D(n2164), .SI(n1338), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4502), .Q(\regfile[9][19] ), .QN(n1337) );
  SDFFNSRXL \regfile_reg[9][18]  ( .D(n2162), .SI(n1339), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4502), .Q(\regfile[9][18] ), .QN(n1338) );
  SDFFNSRXL \regfile_reg[9][17]  ( .D(n2160), .SI(n1340), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4502), .Q(\regfile[9][17] ), .QN(n1339) );
  SDFFNSRXL \regfile_reg[9][16]  ( .D(n2158), .SI(n1341), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4502), .Q(\regfile[9][16] ), .QN(n1340) );
  SDFFNSRXL \regfile_reg[9][15]  ( .D(n2156), .SI(n1342), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4502), .Q(\regfile[9][15] ), .QN(n1341) );
  SDFFNSRXL \regfile_reg[9][14]  ( .D(n2154), .SI(n1343), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4502), .Q(\regfile[9][14] ), .QN(n1342) );
  SDFFNSRXL \regfile_reg[9][13]  ( .D(n2152), .SI(n1344), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4503), .Q(\regfile[9][13] ), .QN(n1343) );
  SDFFNSRXL \regfile_reg[9][12]  ( .D(n2150), .SI(n1345), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4503), .Q(\regfile[9][12] ), .QN(n1344) );
  SDFFNSRXL \regfile_reg[9][11]  ( .D(n2148), .SI(n1346), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4503), .Q(\regfile[9][11] ), .QN(n1345) );
  SDFFNSRXL \regfile_reg[9][10]  ( .D(n2146), .SI(n1347), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4503), .Q(\regfile[9][10] ), .QN(n1346) );
  SDFFNSRXL \regfile_reg[9][9]  ( .D(n2144), .SI(n1348), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4503), .Q(\regfile[9][9] ), .QN(n1347) );
  SDFFNSRXL \regfile_reg[9][8]  ( .D(n2142), .SI(n1349), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4503), .Q(\regfile[9][8] ), .QN(n1348) );
  SDFFNSRXL \regfile_reg[9][7]  ( .D(n2140), .SI(n1350), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4503), .Q(\regfile[9][7] ), .QN(n1349) );
  SDFFNSRXL \regfile_reg[9][6]  ( .D(n2138), .SI(n1351), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4503), .Q(\regfile[9][6] ), .QN(n1350) );
  SDFFNSRXL \regfile_reg[9][5]  ( .D(n2136), .SI(n1352), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4503), .Q(\regfile[9][5] ), .QN(n1351) );
  SDFFNSRXL \regfile_reg[9][4]  ( .D(n2134), .SI(n1353), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4503), .Q(\regfile[9][4] ), .QN(n1352) );
  SDFFNSRXL \regfile_reg[9][3]  ( .D(n2132), .SI(n1354), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4503), .Q(\regfile[9][3] ), .QN(n1353) );
  SDFFNSRXL \regfile_reg[9][2]  ( .D(n2130), .SI(n1355), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4503), .Q(\regfile[9][2] ), .QN(n1354) );
  SDFFNSRXL \regfile_reg[9][1]  ( .D(n2128), .SI(n1356), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4503), .Q(\regfile[9][1] ), .QN(n1355) );
  SDFFNSRXL \regfile_reg[9][0]  ( .D(n2126), .SI(n1357), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4503), .Q(\regfile[9][0] ), .QN(n1356) );
  SDFFNSRXL \regfile_reg[5][31]  ( .D(n1932), .SI(n1454), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4509), .Q(\regfile[5][31] ), .QN(n1453) );
  SDFFNSRXL \regfile_reg[5][30]  ( .D(n1930), .SI(n1455), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4509), .Q(\regfile[5][30] ), .QN(n1454) );
  SDFFNSRXL \regfile_reg[5][29]  ( .D(n1928), .SI(n1456), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4509), .Q(\regfile[5][29] ), .QN(n1455) );
  SDFFNSRXL \regfile_reg[5][28]  ( .D(n1926), .SI(n1457), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4509), .Q(\regfile[5][28] ), .QN(n1456) );
  SDFFNSRXL \regfile_reg[5][27]  ( .D(n1924), .SI(n1458), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4509), .Q(\regfile[5][27] ), .QN(n1457) );
  SDFFNSRXL \regfile_reg[5][26]  ( .D(n1922), .SI(n1459), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4509), .Q(\regfile[5][26] ), .QN(n1458) );
  SDFFNSRXL \regfile_reg[5][25]  ( .D(n1920), .SI(n1460), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4509), .Q(\regfile[5][25] ), .QN(n1459) );
  SDFFNSRXL \regfile_reg[5][24]  ( .D(n1918), .SI(n1461), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4509), .Q(\regfile[5][24] ), .QN(n1460) );
  SDFFNSRXL \regfile_reg[5][23]  ( .D(n1916), .SI(n1462), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4509), .Q(\regfile[5][23] ), .QN(n1461) );
  SDFFNSRXL \regfile_reg[5][22]  ( .D(n1914), .SI(n1463), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4509), .Q(\regfile[5][22] ), .QN(n1462) );
  SDFFNSRXL \regfile_reg[5][21]  ( .D(n1912), .SI(n1464), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4509), .Q(\regfile[5][21] ), .QN(n1463) );
  SDFFNSRXL \regfile_reg[5][20]  ( .D(n1910), .SI(n1465), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4509), .Q(\regfile[5][20] ), .QN(n1464) );
  SDFFNSRXL \regfile_reg[5][19]  ( .D(n1908), .SI(n1466), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4509), .Q(\regfile[5][19] ), .QN(n1465) );
  SDFFNSRXL \regfile_reg[5][18]  ( .D(n1906), .SI(n1467), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4509), .Q(\regfile[5][18] ), .QN(n1466) );
  SDFFNSRXL \regfile_reg[5][17]  ( .D(n1904), .SI(n1468), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4509), .Q(\regfile[5][17] ), .QN(n1467) );
  SDFFNSRXL \regfile_reg[5][16]  ( .D(n1902), .SI(n1469), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4509), .Q(\regfile[5][16] ), .QN(n1468) );
  SDFFNSRXL \regfile_reg[5][15]  ( .D(n1900), .SI(n1470), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4510), .Q(\regfile[5][15] ), .QN(n1469) );
  SDFFNSRXL \regfile_reg[5][14]  ( .D(n1898), .SI(n1471), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4510), .Q(\regfile[5][14] ), .QN(n1470) );
  SDFFNSRXL \regfile_reg[5][13]  ( .D(n1896), .SI(n1472), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4510), .Q(\regfile[5][13] ), .QN(n1471) );
  SDFFNSRXL \regfile_reg[5][12]  ( .D(n1894), .SI(n1473), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4510), .Q(\regfile[5][12] ), .QN(n1472) );
  SDFFNSRXL \regfile_reg[5][11]  ( .D(n1892), .SI(n1474), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4510), .Q(\regfile[5][11] ), .QN(n1473) );
  SDFFNSRXL \regfile_reg[5][10]  ( .D(n1890), .SI(n1475), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4510), .Q(\regfile[5][10] ), .QN(n1474) );
  SDFFNSRXL \regfile_reg[5][9]  ( .D(n1888), .SI(n1476), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4510), .Q(\regfile[5][9] ), .QN(n1475) );
  SDFFNSRXL \regfile_reg[5][8]  ( .D(n1886), .SI(n1477), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4510), .Q(\regfile[5][8] ), .QN(n1476) );
  SDFFNSRXL \regfile_reg[5][7]  ( .D(n1884), .SI(n1478), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4510), .Q(\regfile[5][7] ), .QN(n1477) );
  SDFFNSRXL \regfile_reg[5][6]  ( .D(n1882), .SI(n1479), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4510), .Q(\regfile[5][6] ), .QN(n1478) );
  SDFFNSRXL \regfile_reg[5][5]  ( .D(n1880), .SI(n1480), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4510), .Q(\regfile[5][5] ), .QN(n1479) );
  SDFFNSRXL \regfile_reg[5][4]  ( .D(n1878), .SI(n1481), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4510), .Q(\regfile[5][4] ), .QN(n1480) );
  SDFFNSRXL \regfile_reg[5][3]  ( .D(n1876), .SI(n1482), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4510), .Q(\regfile[5][3] ), .QN(n1481) );
  SDFFNSRXL \regfile_reg[5][2]  ( .D(n1874), .SI(n1483), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4510), .Q(\regfile[5][2] ), .QN(n1482) );
  SDFFNSRXL \regfile_reg[5][1]  ( .D(n1872), .SI(n1484), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4510), .Q(\regfile[5][1] ), .QN(n1483) );
  SDFFNSRXL \regfile_reg[5][0]  ( .D(n1870), .SI(n1485), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4510), .Q(\regfile[5][0] ), .QN(n1484) );
  SDFFNSRXL \regfile_reg[28][31]  ( .D(n3404), .SI(n718), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4468), .Q(\regfile[28][31] ), .QN(n717) );
  SDFFNSRXL \regfile_reg[28][30]  ( .D(n3402), .SI(n719), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4468), .Q(\regfile[28][30] ), .QN(n718) );
  SDFFNSRXL \regfile_reg[28][29]  ( .D(n3400), .SI(n720), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4468), .Q(\regfile[28][29] ), .QN(n719) );
  SDFFNSRXL \regfile_reg[28][28]  ( .D(n3398), .SI(n721), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4468), .Q(\regfile[28][28] ), .QN(n720) );
  SDFFNSRXL \regfile_reg[28][27]  ( .D(n3396), .SI(n722), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4468), .Q(\regfile[28][27] ), .QN(n721) );
  SDFFNSRXL \regfile_reg[28][26]  ( .D(n3394), .SI(n723), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4468), .Q(\regfile[28][26] ), .QN(n722) );
  SDFFNSRXL \regfile_reg[28][25]  ( .D(n3392), .SI(n724), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4468), .Q(\regfile[28][25] ), .QN(n723) );
  SDFFNSRXL \regfile_reg[28][24]  ( .D(n3390), .SI(n725), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4468), .Q(\regfile[28][24] ), .QN(n724) );
  SDFFNSRXL \regfile_reg[28][23]  ( .D(n3388), .SI(n726), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4468), .Q(\regfile[28][23] ), .QN(n725) );
  SDFFNSRXL \regfile_reg[28][22]  ( .D(n3386), .SI(n727), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4468), .Q(\regfile[28][22] ), .QN(n726) );
  SDFFNSRXL \regfile_reg[28][21]  ( .D(n3384), .SI(n728), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4468), .Q(\regfile[28][21] ), .QN(n727) );
  SDFFNSRXL \regfile_reg[28][20]  ( .D(n3382), .SI(n729), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4468), .Q(\regfile[28][20] ), .QN(n728) );
  SDFFNSRXL \regfile_reg[28][19]  ( .D(n3380), .SI(n730), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4468), .Q(\regfile[28][19] ), .QN(n729) );
  SDFFNSRXL \regfile_reg[28][18]  ( .D(n3378), .SI(n731), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4468), .Q(\regfile[28][18] ), .QN(n730) );
  SDFFNSRXL \regfile_reg[28][17]  ( .D(n3376), .SI(n732), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4469), .Q(\regfile[28][17] ), .QN(n731) );
  SDFFNSRXL \regfile_reg[28][16]  ( .D(n3374), .SI(n733), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4469), .Q(\regfile[28][16] ), .QN(n732) );
  SDFFNSRXL \regfile_reg[28][15]  ( .D(n3372), .SI(n734), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4469), .Q(\regfile[28][15] ), .QN(n733) );
  SDFFNSRXL \regfile_reg[28][14]  ( .D(n3370), .SI(n735), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4469), .Q(\regfile[28][14] ), .QN(n734) );
  SDFFNSRXL \regfile_reg[28][13]  ( .D(n3368), .SI(n736), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4469), .Q(\regfile[28][13] ), .QN(n735) );
  SDFFNSRXL \regfile_reg[28][12]  ( .D(n3366), .SI(n737), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4469), .Q(\regfile[28][12] ), .QN(n736) );
  SDFFNSRXL \regfile_reg[28][11]  ( .D(n3364), .SI(n738), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4469), .Q(\regfile[28][11] ), .QN(n737) );
  SDFFNSRXL \regfile_reg[28][10]  ( .D(n3362), .SI(n739), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4469), .Q(\regfile[28][10] ), .QN(n738) );
  SDFFNSRXL \regfile_reg[28][9]  ( .D(n3360), .SI(n740), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4469), .Q(\regfile[28][9] ), .QN(n739) );
  SDFFNSRXL \regfile_reg[28][8]  ( .D(n3358), .SI(n741), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4469), .Q(\regfile[28][8] ), .QN(n740) );
  SDFFNSRXL \regfile_reg[28][7]  ( .D(n3356), .SI(n742), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4469), .Q(\regfile[28][7] ), .QN(n741) );
  SDFFNSRXL \regfile_reg[28][6]  ( .D(n3354), .SI(n743), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4469), .Q(\regfile[28][6] ), .QN(n742) );
  SDFFNSRXL \regfile_reg[28][5]  ( .D(n3352), .SI(n744), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4469), .Q(\regfile[28][5] ), .QN(n743) );
  SDFFNSRXL \regfile_reg[28][4]  ( .D(n3350), .SI(n745), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4469), .Q(\regfile[28][4] ), .QN(n744) );
  SDFFNSRXL \regfile_reg[28][3]  ( .D(n3348), .SI(n746), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4469), .Q(\regfile[28][3] ), .QN(n745) );
  SDFFNSRXL \regfile_reg[28][2]  ( .D(n3346), .SI(n747), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4469), .Q(\regfile[28][2] ), .QN(n746) );
  SDFFNSRXL \regfile_reg[28][1]  ( .D(n3344), .SI(n748), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4469), .Q(\regfile[28][1] ), .QN(n747) );
  SDFFNSRXL \regfile_reg[28][0]  ( .D(n3342), .SI(n749), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4469), .Q(\regfile[28][0] ), .QN(n748) );
  SDFFNSRXL \regfile_reg[24][31]  ( .D(n3148), .SI(n846), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4475), .Q(\regfile[24][31] ), .QN(n845) );
  SDFFNSRXL \regfile_reg[24][30]  ( .D(n3146), .SI(n847), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4475), .Q(\regfile[24][30] ), .QN(n846) );
  SDFFNSRXL \regfile_reg[24][29]  ( .D(n3144), .SI(n848), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4475), .Q(\regfile[24][29] ), .QN(n847) );
  SDFFNSRXL \regfile_reg[24][28]  ( .D(n3142), .SI(n849), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4475), .Q(\regfile[24][28] ), .QN(n848) );
  SDFFNSRXL \regfile_reg[24][27]  ( .D(n3140), .SI(n850), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4475), .Q(\regfile[24][27] ), .QN(n849) );
  SDFFNSRXL \regfile_reg[24][26]  ( .D(n3138), .SI(n851), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4475), .Q(\regfile[24][26] ), .QN(n850) );
  SDFFNSRXL \regfile_reg[24][25]  ( .D(n3136), .SI(n852), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4475), .Q(\regfile[24][25] ), .QN(n851) );
  SDFFNSRXL \regfile_reg[24][24]  ( .D(n3134), .SI(n853), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4475), .Q(\regfile[24][24] ), .QN(n852) );
  SDFFNSRXL \regfile_reg[24][23]  ( .D(n3132), .SI(n854), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4475), .Q(\regfile[24][23] ), .QN(n853) );
  SDFFNSRXL \regfile_reg[24][22]  ( .D(n3130), .SI(n855), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4475), .Q(\regfile[24][22] ), .QN(n854) );
  SDFFNSRXL \regfile_reg[24][21]  ( .D(n3128), .SI(n856), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4475), .Q(\regfile[24][21] ), .QN(n855) );
  SDFFNSRXL \regfile_reg[24][20]  ( .D(n3126), .SI(n857), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4475), .Q(\regfile[24][20] ), .QN(n856) );
  SDFFNSRXL \regfile_reg[24][19]  ( .D(n3124), .SI(n858), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4476), .Q(\regfile[24][19] ), .QN(n857) );
  SDFFNSRXL \regfile_reg[24][18]  ( .D(n3122), .SI(n859), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4476), .Q(\regfile[24][18] ), .QN(n858) );
  SDFFNSRXL \regfile_reg[24][17]  ( .D(n3120), .SI(n860), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4476), .Q(\regfile[24][17] ), .QN(n859) );
  SDFFNSRXL \regfile_reg[24][16]  ( .D(n3118), .SI(n861), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4476), .Q(\regfile[24][16] ), .QN(n860) );
  SDFFNSRXL \regfile_reg[24][15]  ( .D(n3116), .SI(n862), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4476), .Q(\regfile[24][15] ), .QN(n861) );
  SDFFNSRXL \regfile_reg[24][14]  ( .D(n3114), .SI(n863), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4476), .Q(\regfile[24][14] ), .QN(n862) );
  SDFFNSRXL \regfile_reg[24][13]  ( .D(n3112), .SI(n864), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4476), .Q(\regfile[24][13] ), .QN(n863) );
  SDFFNSRXL \regfile_reg[24][12]  ( .D(n3110), .SI(n865), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4476), .Q(\regfile[24][12] ), .QN(n864) );
  SDFFNSRXL \regfile_reg[24][11]  ( .D(n3108), .SI(n866), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4476), .Q(\regfile[24][11] ), .QN(n865) );
  SDFFNSRXL \regfile_reg[24][10]  ( .D(n3106), .SI(n867), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4476), .Q(\regfile[24][10] ), .QN(n866) );
  SDFFNSRXL \regfile_reg[24][9]  ( .D(n3104), .SI(n868), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4476), .Q(\regfile[24][9] ), .QN(n867) );
  SDFFNSRXL \regfile_reg[24][8]  ( .D(n3102), .SI(n869), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4476), .Q(\regfile[24][8] ), .QN(n868) );
  SDFFNSRXL \regfile_reg[24][7]  ( .D(n3100), .SI(n870), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4476), .Q(\regfile[24][7] ), .QN(n869) );
  SDFFNSRXL \regfile_reg[24][6]  ( .D(n3098), .SI(n871), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4476), .Q(\regfile[24][6] ), .QN(n870) );
  SDFFNSRXL \regfile_reg[24][5]  ( .D(n3096), .SI(n872), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4476), .Q(\regfile[24][5] ), .QN(n871) );
  SDFFNSRXL \regfile_reg[24][4]  ( .D(n3094), .SI(n873), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4476), .Q(\regfile[24][4] ), .QN(n872) );
  SDFFNSRXL \regfile_reg[24][3]  ( .D(n3092), .SI(n874), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4476), .Q(\regfile[24][3] ), .QN(n873) );
  SDFFNSRXL \regfile_reg[24][2]  ( .D(n3090), .SI(n875), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4476), .Q(\regfile[24][2] ), .QN(n874) );
  SDFFNSRXL \regfile_reg[24][1]  ( .D(n3088), .SI(n876), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4477), .Q(\regfile[24][1] ), .QN(n875) );
  SDFFNSRXL \regfile_reg[24][0]  ( .D(n3086), .SI(n877), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4477), .Q(\regfile[24][0] ), .QN(n876) );
  SDFFNSRXL \regfile_reg[20][31]  ( .D(n2892), .SI(n974), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4482), .Q(\regfile[20][31] ), .QN(n973) );
  SDFFNSRXL \regfile_reg[20][30]  ( .D(n2890), .SI(n975), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4482), .Q(\regfile[20][30] ), .QN(n974) );
  SDFFNSRXL \regfile_reg[20][29]  ( .D(n2888), .SI(n976), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4482), .Q(\regfile[20][29] ), .QN(n975) );
  SDFFNSRXL \regfile_reg[20][28]  ( .D(n2886), .SI(n977), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4482), .Q(\regfile[20][28] ), .QN(n976) );
  SDFFNSRXL \regfile_reg[20][27]  ( .D(n2884), .SI(n978), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4482), .Q(\regfile[20][27] ), .QN(n977) );
  SDFFNSRXL \regfile_reg[20][26]  ( .D(n2882), .SI(n979), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4482), .Q(\regfile[20][26] ), .QN(n978) );
  SDFFNSRXL \regfile_reg[20][25]  ( .D(n2880), .SI(n980), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4482), .Q(\regfile[20][25] ), .QN(n979) );
  SDFFNSRXL \regfile_reg[20][24]  ( .D(n2878), .SI(n981), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4482), .Q(\regfile[20][24] ), .QN(n980) );
  SDFFNSRXL \regfile_reg[20][23]  ( .D(n2876), .SI(n982), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4482), .Q(\regfile[20][23] ), .QN(n981) );
  SDFFNSRXL \regfile_reg[20][22]  ( .D(n2874), .SI(n983), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4482), .Q(\regfile[20][22] ), .QN(n982) );
  SDFFNSRXL \regfile_reg[20][21]  ( .D(n2872), .SI(n984), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4483), .Q(\regfile[20][21] ), .QN(n983) );
  SDFFNSRXL \regfile_reg[20][20]  ( .D(n2870), .SI(n985), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4483), .Q(\regfile[20][20] ), .QN(n984) );
  SDFFNSRXL \regfile_reg[20][19]  ( .D(n2868), .SI(n986), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4483), .Q(\regfile[20][19] ), .QN(n985) );
  SDFFNSRXL \regfile_reg[20][18]  ( .D(n2866), .SI(n987), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4483), .Q(\regfile[20][18] ), .QN(n986) );
  SDFFNSRXL \regfile_reg[20][17]  ( .D(n2864), .SI(n988), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4483), .Q(\regfile[20][17] ), .QN(n987) );
  SDFFNSRXL \regfile_reg[20][16]  ( .D(n2862), .SI(n989), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4483), .Q(\regfile[20][16] ), .QN(n988) );
  SDFFNSRXL \regfile_reg[20][15]  ( .D(n2860), .SI(n990), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4483), .Q(\regfile[20][15] ), .QN(n989) );
  SDFFNSRXL \regfile_reg[20][14]  ( .D(n2858), .SI(n991), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4483), .Q(\regfile[20][14] ), .QN(n990) );
  SDFFNSRXL \regfile_reg[20][13]  ( .D(n2856), .SI(n992), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4483), .Q(\regfile[20][13] ), .QN(n991) );
  SDFFNSRXL \regfile_reg[20][12]  ( .D(n2854), .SI(n993), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4483), .Q(\regfile[20][12] ), .QN(n992) );
  SDFFNSRXL \regfile_reg[20][11]  ( .D(n2852), .SI(n994), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4483), .Q(\regfile[20][11] ), .QN(n993) );
  SDFFNSRXL \regfile_reg[20][10]  ( .D(n2850), .SI(n995), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4483), .Q(\regfile[20][10] ), .QN(n994) );
  SDFFNSRXL \regfile_reg[20][9]  ( .D(n2848), .SI(n996), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4483), .Q(\regfile[20][9] ), .QN(n995) );
  SDFFNSRXL \regfile_reg[20][8]  ( .D(n2846), .SI(n997), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4483), .Q(\regfile[20][8] ), .QN(n996) );
  SDFFNSRXL \regfile_reg[20][7]  ( .D(n2844), .SI(n998), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4483), .Q(\regfile[20][7] ), .QN(n997) );
  SDFFNSRXL \regfile_reg[20][6]  ( .D(n2842), .SI(n999), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4483), .Q(\regfile[20][6] ), .QN(n998) );
  SDFFNSRXL \regfile_reg[20][5]  ( .D(n2840), .SI(n1000), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4483), .Q(\regfile[20][5] ), .QN(n999) );
  SDFFNSRXL \regfile_reg[20][4]  ( .D(n2838), .SI(n1001), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4483), .Q(\regfile[20][4] ), .QN(n1000) );
  SDFFNSRXL \regfile_reg[20][3]  ( .D(n2836), .SI(n1002), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4484), .Q(\regfile[20][3] ), .QN(n1001) );
  SDFFNSRXL \regfile_reg[20][2]  ( .D(n2834), .SI(n1003), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4484), .Q(\regfile[20][2] ), .QN(n1002) );
  SDFFNSRXL \regfile_reg[20][1]  ( .D(n2832), .SI(n1004), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4484), .Q(\regfile[20][1] ), .QN(n1003) );
  SDFFNSRXL \regfile_reg[20][0]  ( .D(n2830), .SI(n1005), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4484), .Q(\regfile[20][0] ), .QN(n1004) );
  SDFFNSRXL \regfile_reg[16][31]  ( .D(n2636), .SI(n1102), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4489), .Q(\regfile[16][31] ), .QN(n1101) );
  SDFFNSRXL \regfile_reg[16][30]  ( .D(n2634), .SI(n1103), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4489), .Q(\regfile[16][30] ), .QN(n1102) );
  SDFFNSRXL \regfile_reg[16][29]  ( .D(n2632), .SI(n1104), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4489), .Q(\regfile[16][29] ), .QN(n1103) );
  SDFFNSRXL \regfile_reg[16][28]  ( .D(n2630), .SI(n1105), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4489), .Q(\regfile[16][28] ), .QN(n1104) );
  SDFFNSRXL \regfile_reg[16][27]  ( .D(n2628), .SI(n1106), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4489), .Q(\regfile[16][27] ), .QN(n1105) );
  SDFFNSRXL \regfile_reg[16][26]  ( .D(n2626), .SI(n1107), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4489), .Q(\regfile[16][26] ), .QN(n1106) );
  SDFFNSRXL \regfile_reg[16][25]  ( .D(n2624), .SI(n1108), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4489), .Q(\regfile[16][25] ), .QN(n1107) );
  SDFFNSRXL \regfile_reg[16][24]  ( .D(n2622), .SI(n1109), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4489), .Q(\regfile[16][24] ), .QN(n1108) );
  SDFFNSRXL \regfile_reg[16][23]  ( .D(n2620), .SI(n1110), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4490), .Q(\regfile[16][23] ), .QN(n1109) );
  SDFFNSRXL \regfile_reg[16][22]  ( .D(n2618), .SI(n1111), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4490), .Q(\regfile[16][22] ), .QN(n1110) );
  SDFFNSRXL \regfile_reg[16][21]  ( .D(n2616), .SI(n1112), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4490), .Q(\regfile[16][21] ), .QN(n1111) );
  SDFFNSRXL \regfile_reg[16][20]  ( .D(n2614), .SI(n1113), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4490), .Q(\regfile[16][20] ), .QN(n1112) );
  SDFFNSRXL \regfile_reg[16][19]  ( .D(n2612), .SI(n1114), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4490), .Q(\regfile[16][19] ), .QN(n1113) );
  SDFFNSRXL \regfile_reg[16][18]  ( .D(n2610), .SI(n1115), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4490), .Q(\regfile[16][18] ), .QN(n1114) );
  SDFFNSRXL \regfile_reg[16][17]  ( .D(n2608), .SI(n1116), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4490), .Q(\regfile[16][17] ), .QN(n1115) );
  SDFFNSRXL \regfile_reg[16][16]  ( .D(n2606), .SI(n1117), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4490), .Q(\regfile[16][16] ), .QN(n1116) );
  SDFFNSRXL \regfile_reg[16][15]  ( .D(n2604), .SI(n1118), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4490), .Q(\regfile[16][15] ), .QN(n1117) );
  SDFFNSRXL \regfile_reg[16][14]  ( .D(n2602), .SI(n1119), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4490), .Q(\regfile[16][14] ), .QN(n1118) );
  SDFFNSRXL \regfile_reg[16][13]  ( .D(n2600), .SI(n1120), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4490), .Q(\regfile[16][13] ), .QN(n1119) );
  SDFFNSRXL \regfile_reg[16][12]  ( .D(n2598), .SI(n1121), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4490), .Q(\regfile[16][12] ), .QN(n1120) );
  SDFFNSRXL \regfile_reg[16][11]  ( .D(n2596), .SI(n1122), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4490), .Q(\regfile[16][11] ), .QN(n1121) );
  SDFFNSRXL \regfile_reg[16][10]  ( .D(n2594), .SI(n1123), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4490), .Q(\regfile[16][10] ), .QN(n1122) );
  SDFFNSRXL \regfile_reg[16][9]  ( .D(n2592), .SI(n1124), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4490), .Q(\regfile[16][9] ), .QN(n1123) );
  SDFFNSRXL \regfile_reg[16][8]  ( .D(n2590), .SI(n1125), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4490), .Q(\regfile[16][8] ), .QN(n1124) );
  SDFFNSRXL \regfile_reg[16][7]  ( .D(n2588), .SI(n1126), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4490), .Q(\regfile[16][7] ), .QN(n1125) );
  SDFFNSRXL \regfile_reg[16][6]  ( .D(n2586), .SI(n1127), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4490), .Q(\regfile[16][6] ), .QN(n1126) );
  SDFFNSRXL \regfile_reg[16][5]  ( .D(n2584), .SI(n1128), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4491), .Q(\regfile[16][5] ), .QN(n1127) );
  SDFFNSRXL \regfile_reg[16][4]  ( .D(n2582), .SI(n1129), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4491), .Q(\regfile[16][4] ), .QN(n1128) );
  SDFFNSRXL \regfile_reg[16][3]  ( .D(n2580), .SI(n1130), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4491), .Q(\regfile[16][3] ), .QN(n1129) );
  SDFFNSRXL \regfile_reg[16][2]  ( .D(n2578), .SI(n1131), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4491), .Q(\regfile[16][2] ), .QN(n1130) );
  SDFFNSRXL \regfile_reg[16][1]  ( .D(n2576), .SI(n1132), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4491), .Q(\regfile[16][1] ), .QN(n1131) );
  SDFFNSRXL \regfile_reg[16][0]  ( .D(n2574), .SI(n1133), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4491), .Q(\regfile[16][0] ), .QN(n1132) );
  SDFFNSRXL \regfile_reg[12][31]  ( .D(n2380), .SI(n1230), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4496), .Q(\regfile[12][31] ), .QN(n1229) );
  SDFFNSRXL \regfile_reg[12][30]  ( .D(n2378), .SI(n1231), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4496), .Q(\regfile[12][30] ), .QN(n1230) );
  SDFFNSRXL \regfile_reg[12][29]  ( .D(n2376), .SI(n1232), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4496), .Q(\regfile[12][29] ), .QN(n1231) );
  SDFFNSRXL \regfile_reg[12][28]  ( .D(n2374), .SI(n1233), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4496), .Q(\regfile[12][28] ), .QN(n1232) );
  SDFFNSRXL \regfile_reg[12][27]  ( .D(n2372), .SI(n1234), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4496), .Q(\regfile[12][27] ), .QN(n1233) );
  SDFFNSRXL \regfile_reg[12][26]  ( .D(n2370), .SI(n1235), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4496), .Q(\regfile[12][26] ), .QN(n1234) );
  SDFFNSRXL \regfile_reg[12][25]  ( .D(n2368), .SI(n1236), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4497), .Q(\regfile[12][25] ), .QN(n1235) );
  SDFFNSRXL \regfile_reg[12][24]  ( .D(n2366), .SI(n1237), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4497), .Q(\regfile[12][24] ), .QN(n1236) );
  SDFFNSRXL \regfile_reg[12][23]  ( .D(n2364), .SI(n1238), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4497), .Q(\regfile[12][23] ), .QN(n1237) );
  SDFFNSRXL \regfile_reg[12][22]  ( .D(n2362), .SI(n1239), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4497), .Q(\regfile[12][22] ), .QN(n1238) );
  SDFFNSRXL \regfile_reg[12][21]  ( .D(n2360), .SI(n1240), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4497), .Q(\regfile[12][21] ), .QN(n1239) );
  SDFFNSRXL \regfile_reg[12][20]  ( .D(n2358), .SI(n1241), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4497), .Q(\regfile[12][20] ), .QN(n1240) );
  SDFFNSRXL \regfile_reg[12][19]  ( .D(n2356), .SI(n1242), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4497), .Q(\regfile[12][19] ), .QN(n1241) );
  SDFFNSRXL \regfile_reg[12][18]  ( .D(n2354), .SI(n1243), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4497), .Q(\regfile[12][18] ), .QN(n1242) );
  SDFFNSRXL \regfile_reg[12][17]  ( .D(n2352), .SI(n1244), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4497), .Q(\regfile[12][17] ), .QN(n1243) );
  SDFFNSRXL \regfile_reg[12][16]  ( .D(n2350), .SI(n1245), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4497), .Q(\regfile[12][16] ), .QN(n1244) );
  SDFFNSRXL \regfile_reg[12][15]  ( .D(n2348), .SI(n1246), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4497), .Q(\regfile[12][15] ), .QN(n1245) );
  SDFFNSRXL \regfile_reg[12][14]  ( .D(n2346), .SI(n1247), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4497), .Q(\regfile[12][14] ), .QN(n1246) );
  SDFFNSRXL \regfile_reg[12][13]  ( .D(n2344), .SI(n1248), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4497), .Q(\regfile[12][13] ), .QN(n1247) );
  SDFFNSRXL \regfile_reg[12][12]  ( .D(n2342), .SI(n1249), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4497), .Q(\regfile[12][12] ), .QN(n1248) );
  SDFFNSRXL \regfile_reg[12][11]  ( .D(n2340), .SI(n1250), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4497), .Q(\regfile[12][11] ), .QN(n1249) );
  SDFFNSRXL \regfile_reg[12][10]  ( .D(n2338), .SI(n1251), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4497), .Q(\regfile[12][10] ), .QN(n1250) );
  SDFFNSRXL \regfile_reg[12][9]  ( .D(n2336), .SI(n1252), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4497), .Q(\regfile[12][9] ), .QN(n1251) );
  SDFFNSRXL \regfile_reg[12][8]  ( .D(n2334), .SI(n1253), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4497), .Q(\regfile[12][8] ), .QN(n1252) );
  SDFFNSRXL \regfile_reg[12][7]  ( .D(n2332), .SI(n1254), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4498), .Q(\regfile[12][7] ), .QN(n1253) );
  SDFFNSRXL \regfile_reg[12][6]  ( .D(n2330), .SI(n1255), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4498), .Q(\regfile[12][6] ), .QN(n1254) );
  SDFFNSRXL \regfile_reg[12][5]  ( .D(n2328), .SI(n1256), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4498), .Q(\regfile[12][5] ), .QN(n1255) );
  SDFFNSRXL \regfile_reg[12][4]  ( .D(n2326), .SI(n1257), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4498), .Q(\regfile[12][4] ), .QN(n1256) );
  SDFFNSRXL \regfile_reg[12][3]  ( .D(n2324), .SI(n1258), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4498), .Q(\regfile[12][3] ), .QN(n1257) );
  SDFFNSRXL \regfile_reg[12][2]  ( .D(n2322), .SI(n1259), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4498), .Q(\regfile[12][2] ), .QN(n1258) );
  SDFFNSRXL \regfile_reg[12][1]  ( .D(n2320), .SI(n1260), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4498), .Q(\regfile[12][1] ), .QN(n1259) );
  SDFFNSRXL \regfile_reg[12][0]  ( .D(n2318), .SI(n1261), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4498), .Q(\regfile[12][0] ), .QN(n1260) );
  SDFFNSRXL \regfile_reg[8][31]  ( .D(n2124), .SI(n1358), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4503), .Q(\regfile[8][31] ), .QN(n1357) );
  SDFFNSRXL \regfile_reg[8][30]  ( .D(n2122), .SI(n1359), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4503), .Q(\regfile[8][30] ), .QN(n1358) );
  SDFFNSRXL \regfile_reg[8][29]  ( .D(n2120), .SI(n1360), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4503), .Q(\regfile[8][29] ), .QN(n1359) );
  SDFFNSRXL \regfile_reg[8][28]  ( .D(n2118), .SI(n1361), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4503), .Q(\regfile[8][28] ), .QN(n1360) );
  SDFFNSRXL \regfile_reg[8][27]  ( .D(n2116), .SI(n1362), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4504), .Q(\regfile[8][27] ), .QN(n1361) );
  SDFFNSRXL \regfile_reg[8][26]  ( .D(n2114), .SI(n1363), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4504), .Q(\regfile[8][26] ), .QN(n1362) );
  SDFFNSRXL \regfile_reg[8][25]  ( .D(n2112), .SI(n1364), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4504), .Q(\regfile[8][25] ), .QN(n1363) );
  SDFFNSRXL \regfile_reg[8][24]  ( .D(n2110), .SI(n1365), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4504), .Q(\regfile[8][24] ), .QN(n1364) );
  SDFFNSRXL \regfile_reg[8][23]  ( .D(n2108), .SI(n1366), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4504), .Q(\regfile[8][23] ), .QN(n1365) );
  SDFFNSRXL \regfile_reg[8][22]  ( .D(n2106), .SI(n1367), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4504), .Q(\regfile[8][22] ), .QN(n1366) );
  SDFFNSRXL \regfile_reg[8][21]  ( .D(n2104), .SI(n1368), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4504), .Q(\regfile[8][21] ), .QN(n1367) );
  SDFFNSRXL \regfile_reg[8][20]  ( .D(n2102), .SI(n1369), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4504), .Q(\regfile[8][20] ), .QN(n1368) );
  SDFFNSRXL \regfile_reg[8][19]  ( .D(n2100), .SI(n1370), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4504), .Q(\regfile[8][19] ), .QN(n1369) );
  SDFFNSRXL \regfile_reg[8][18]  ( .D(n2098), .SI(n1371), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4504), .Q(\regfile[8][18] ), .QN(n1370) );
  SDFFNSRXL \regfile_reg[8][17]  ( .D(n2096), .SI(n1372), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4504), .Q(\regfile[8][17] ), .QN(n1371) );
  SDFFNSRXL \regfile_reg[8][16]  ( .D(n2094), .SI(n1373), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4504), .Q(\regfile[8][16] ), .QN(n1372) );
  SDFFNSRXL \regfile_reg[8][15]  ( .D(n2092), .SI(n1374), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4504), .Q(\regfile[8][15] ), .QN(n1373) );
  SDFFNSRXL \regfile_reg[8][14]  ( .D(n2090), .SI(n1375), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4504), .Q(\regfile[8][14] ), .QN(n1374) );
  SDFFNSRXL \regfile_reg[8][13]  ( .D(n2088), .SI(n1376), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4504), .Q(\regfile[8][13] ), .QN(n1375) );
  SDFFNSRXL \regfile_reg[8][12]  ( .D(n2086), .SI(n1377), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4504), .Q(\regfile[8][12] ), .QN(n1376) );
  SDFFNSRXL \regfile_reg[8][11]  ( .D(n2084), .SI(n1378), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4504), .Q(\regfile[8][11] ), .QN(n1377) );
  SDFFNSRXL \regfile_reg[8][10]  ( .D(n2082), .SI(n1379), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4504), .Q(\regfile[8][10] ), .QN(n1378) );
  SDFFNSRXL \regfile_reg[8][9]  ( .D(n2080), .SI(n1380), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4505), .Q(\regfile[8][9] ), .QN(n1379) );
  SDFFNSRXL \regfile_reg[8][8]  ( .D(n2078), .SI(n1381), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4505), .Q(\regfile[8][8] ), .QN(n1380) );
  SDFFNSRXL \regfile_reg[8][7]  ( .D(n2076), .SI(n1382), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4505), .Q(\regfile[8][7] ), .QN(n1381) );
  SDFFNSRXL \regfile_reg[8][6]  ( .D(n2074), .SI(n1383), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4505), .Q(\regfile[8][6] ), .QN(n1382) );
  SDFFNSRXL \regfile_reg[8][5]  ( .D(n2072), .SI(n1384), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4505), .Q(\regfile[8][5] ), .QN(n1383) );
  SDFFNSRXL \regfile_reg[8][4]  ( .D(n2070), .SI(n1385), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4505), .Q(\regfile[8][4] ), .QN(n1384) );
  SDFFNSRXL \regfile_reg[8][3]  ( .D(n2068), .SI(n1386), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4505), .Q(\regfile[8][3] ), .QN(n1385) );
  SDFFNSRXL \regfile_reg[8][2]  ( .D(n2066), .SI(n1387), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4505), .Q(\regfile[8][2] ), .QN(n1386) );
  SDFFNSRXL \regfile_reg[8][1]  ( .D(n2064), .SI(n1388), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4505), .Q(\regfile[8][1] ), .QN(n1387) );
  SDFFNSRXL \regfile_reg[8][0]  ( .D(n2062), .SI(n1389), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4505), .Q(\regfile[8][0] ), .QN(n1388) );
  SDFFNSRXL \regfile_reg[4][31]  ( .D(n1868), .SI(n1486), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4510), .Q(\regfile[4][31] ), .QN(n1485) );
  SDFFNSRXL \regfile_reg[4][30]  ( .D(n1866), .SI(n1487), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4510), .Q(\regfile[4][30] ), .QN(n1486) );
  SDFFNSRXL \regfile_reg[4][29]  ( .D(n1864), .SI(n1488), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4511), .Q(\regfile[4][29] ), .QN(n1487) );
  SDFFNSRXL \regfile_reg[4][28]  ( .D(n1862), .SI(n1489), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4511), .Q(\regfile[4][28] ), .QN(n1488) );
  SDFFNSRXL \regfile_reg[4][27]  ( .D(n1860), .SI(n1490), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4511), .Q(\regfile[4][27] ), .QN(n1489) );
  SDFFNSRXL \regfile_reg[4][26]  ( .D(n1858), .SI(n1491), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4511), .Q(\regfile[4][26] ), .QN(n1490) );
  SDFFNSRXL \regfile_reg[4][25]  ( .D(n1856), .SI(n1492), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4511), .Q(\regfile[4][25] ), .QN(n1491) );
  SDFFNSRXL \regfile_reg[4][24]  ( .D(n1854), .SI(n1493), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4511), .Q(\regfile[4][24] ), .QN(n1492) );
  SDFFNSRXL \regfile_reg[4][23]  ( .D(n1852), .SI(n1494), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4511), .Q(\regfile[4][23] ), .QN(n1493) );
  SDFFNSRXL \regfile_reg[4][22]  ( .D(n1850), .SI(n1495), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4511), .Q(\regfile[4][22] ), .QN(n1494) );
  SDFFNSRXL \regfile_reg[4][21]  ( .D(n1848), .SI(n1496), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4511), .Q(\regfile[4][21] ), .QN(n1495) );
  SDFFNSRXL \regfile_reg[4][20]  ( .D(n1846), .SI(n1497), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4511), .Q(\regfile[4][20] ), .QN(n1496) );
  SDFFNSRXL \regfile_reg[4][19]  ( .D(n1844), .SI(n1498), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4511), .Q(\regfile[4][19] ), .QN(n1497) );
  SDFFNSRXL \regfile_reg[4][18]  ( .D(n1842), .SI(n1499), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4511), .Q(\regfile[4][18] ), .QN(n1498) );
  SDFFNSRXL \regfile_reg[4][17]  ( .D(n1840), .SI(n1500), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4511), .Q(\regfile[4][17] ), .QN(n1499) );
  SDFFNSRXL \regfile_reg[4][16]  ( .D(n1838), .SI(n1501), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4511), .Q(\regfile[4][16] ), .QN(n1500) );
  SDFFNSRXL \regfile_reg[4][15]  ( .D(n1836), .SI(n1502), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4511), .Q(\regfile[4][15] ), .QN(n1501) );
  SDFFNSRXL \regfile_reg[4][14]  ( .D(n1834), .SI(n1503), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4511), .Q(\regfile[4][14] ), .QN(n1502) );
  SDFFNSRXL \regfile_reg[4][13]  ( .D(n1832), .SI(n1504), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4511), .Q(\regfile[4][13] ), .QN(n1503) );
  SDFFNSRXL \regfile_reg[4][12]  ( .D(n1830), .SI(n1505), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4511), .Q(\regfile[4][12] ), .QN(n1504) );
  SDFFNSRXL \regfile_reg[4][11]  ( .D(n1828), .SI(n1506), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4512), .Q(\regfile[4][11] ), .QN(n1505) );
  SDFFNSRXL \regfile_reg[4][10]  ( .D(n1826), .SI(n1507), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4512), .Q(\regfile[4][10] ), .QN(n1506) );
  SDFFNSRXL \regfile_reg[4][9]  ( .D(n1824), .SI(n1508), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4512), .Q(\regfile[4][9] ), .QN(n1507) );
  SDFFNSRXL \regfile_reg[4][8]  ( .D(n1822), .SI(n1509), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4512), .Q(\regfile[4][8] ), .QN(n1508) );
  SDFFNSRXL \regfile_reg[4][7]  ( .D(n1820), .SI(n1510), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4512), .Q(\regfile[4][7] ), .QN(n1509) );
  SDFFNSRXL \regfile_reg[4][6]  ( .D(n1818), .SI(n1511), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4512), .Q(\regfile[4][6] ), .QN(n1510) );
  SDFFNSRXL \regfile_reg[4][5]  ( .D(n1816), .SI(n1512), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4512), .Q(\regfile[4][5] ), .QN(n1511) );
  SDFFNSRXL \regfile_reg[4][4]  ( .D(n1814), .SI(n1513), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4512), .Q(\regfile[4][4] ), .QN(n1512) );
  SDFFNSRXL \regfile_reg[4][3]  ( .D(n1812), .SI(n1514), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4512), .Q(\regfile[4][3] ), .QN(n1513) );
  SDFFNSRXL \regfile_reg[4][2]  ( .D(n1810), .SI(n1515), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4512), .Q(\regfile[4][2] ), .QN(n1514) );
  SDFFNSRXL \regfile_reg[4][1]  ( .D(n1808), .SI(n1516), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4512), .Q(\regfile[4][1] ), .QN(n1515) );
  SDFFNSRXL \regfile_reg[4][0]  ( .D(n1806), .SI(n1517), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4512), .Q(\regfile[4][0] ), .QN(n1516) );
  SDFFNSRXL \regfile_reg[30][31]  ( .D(n3532), .SI(n654), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4464), .Q(\regfile[30][31] ), .QN(n653) );
  SDFFNSRXL \regfile_reg[30][30]  ( .D(n3530), .SI(n655), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4464), .Q(\regfile[30][30] ), .QN(n654) );
  SDFFNSRXL \regfile_reg[30][29]  ( .D(n3528), .SI(n656), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4464), .Q(\regfile[30][29] ), .QN(n655) );
  SDFFNSRXL \regfile_reg[30][28]  ( .D(n3526), .SI(n657), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4464), .Q(\regfile[30][28] ), .QN(n656) );
  SDFFNSRXL \regfile_reg[30][27]  ( .D(n3524), .SI(n658), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4464), .Q(\regfile[30][27] ), .QN(n657) );
  SDFFNSRXL \regfile_reg[30][26]  ( .D(n3522), .SI(n659), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4464), .Q(\regfile[30][26] ), .QN(n658) );
  SDFFNSRXL \regfile_reg[30][25]  ( .D(n3520), .SI(n660), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4465), .Q(\regfile[30][25] ), .QN(n659) );
  SDFFNSRXL \regfile_reg[30][24]  ( .D(n3518), .SI(n661), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4465), .Q(\regfile[30][24] ), .QN(n660) );
  SDFFNSRXL \regfile_reg[30][23]  ( .D(n3516), .SI(n662), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4465), .Q(\regfile[30][23] ), .QN(n661) );
  SDFFNSRXL \regfile_reg[30][22]  ( .D(n3514), .SI(n663), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4465), .Q(\regfile[30][22] ), .QN(n662) );
  SDFFNSRXL \regfile_reg[30][21]  ( .D(n3512), .SI(n664), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4465), .Q(\regfile[30][21] ), .QN(n663) );
  SDFFNSRXL \regfile_reg[30][20]  ( .D(n3510), .SI(n665), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4465), .Q(\regfile[30][20] ), .QN(n664) );
  SDFFNSRXL \regfile_reg[30][19]  ( .D(n3508), .SI(n666), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4465), .Q(\regfile[30][19] ), .QN(n665) );
  SDFFNSRXL \regfile_reg[30][18]  ( .D(n3506), .SI(n667), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4465), .Q(\regfile[30][18] ), .QN(n666) );
  SDFFNSRXL \regfile_reg[30][17]  ( .D(n3504), .SI(n668), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4465), .Q(\regfile[30][17] ), .QN(n667) );
  SDFFNSRXL \regfile_reg[30][16]  ( .D(n3502), .SI(n669), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4465), .Q(\regfile[30][16] ), .QN(n668) );
  SDFFNSRXL \regfile_reg[30][15]  ( .D(n3500), .SI(n670), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4465), .Q(\regfile[30][15] ), .QN(n669) );
  SDFFNSRXL \regfile_reg[30][14]  ( .D(n3498), .SI(n671), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4465), .Q(\regfile[30][14] ), .QN(n670) );
  SDFFNSRXL \regfile_reg[30][13]  ( .D(n3496), .SI(n672), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4465), .Q(\regfile[30][13] ), .QN(n671) );
  SDFFNSRXL \regfile_reg[30][12]  ( .D(n3494), .SI(n673), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4465), .Q(\regfile[30][12] ), .QN(n672) );
  SDFFNSRXL \regfile_reg[30][11]  ( .D(n3492), .SI(n674), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4465), .Q(\regfile[30][11] ), .QN(n673) );
  SDFFNSRXL \regfile_reg[30][10]  ( .D(n3490), .SI(n675), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4465), .Q(\regfile[30][10] ), .QN(n674) );
  SDFFNSRXL \regfile_reg[30][9]  ( .D(n3488), .SI(n676), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4465), .Q(\regfile[30][9] ), .QN(n675) );
  SDFFNSRXL \regfile_reg[30][8]  ( .D(n3486), .SI(n677), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4465), .Q(\regfile[30][8] ), .QN(n676) );
  SDFFNSRXL \regfile_reg[30][7]  ( .D(n3484), .SI(n678), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4466), .Q(\regfile[30][7] ), .QN(n677) );
  SDFFNSRXL \regfile_reg[30][6]  ( .D(n3482), .SI(n679), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4466), .Q(\regfile[30][6] ), .QN(n678) );
  SDFFNSRXL \regfile_reg[30][5]  ( .D(n3480), .SI(n680), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4466), .Q(\regfile[30][5] ), .QN(n679) );
  SDFFNSRXL \regfile_reg[30][4]  ( .D(n3478), .SI(n681), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4466), .Q(\regfile[30][4] ), .QN(n680) );
  SDFFNSRXL \regfile_reg[30][3]  ( .D(n3476), .SI(n682), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4466), .Q(\regfile[30][3] ), .QN(n681) );
  SDFFNSRXL \regfile_reg[30][2]  ( .D(n3474), .SI(n683), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4466), .Q(\regfile[30][2] ), .QN(n682) );
  SDFFNSRXL \regfile_reg[30][1]  ( .D(n3472), .SI(n684), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4466), .Q(\regfile[30][1] ), .QN(n683) );
  SDFFNSRXL \regfile_reg[30][0]  ( .D(n3470), .SI(n685), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4466), .Q(\regfile[30][0] ), .QN(n684) );
  SDFFNSRXL \regfile_reg[26][31]  ( .D(n3276), .SI(n782), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4471), .Q(\regfile[26][31] ), .QN(n781) );
  SDFFNSRXL \regfile_reg[26][30]  ( .D(n3274), .SI(n783), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4471), .Q(\regfile[26][30] ), .QN(n782) );
  SDFFNSRXL \regfile_reg[26][29]  ( .D(n3272), .SI(n784), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4471), .Q(\regfile[26][29] ), .QN(n783) );
  SDFFNSRXL \regfile_reg[26][28]  ( .D(n3270), .SI(n785), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4471), .Q(\regfile[26][28] ), .QN(n784) );
  SDFFNSRXL \regfile_reg[26][27]  ( .D(n3268), .SI(n786), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4472), .Q(\regfile[26][27] ), .QN(n785) );
  SDFFNSRXL \regfile_reg[26][26]  ( .D(n3266), .SI(n787), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4472), .Q(\regfile[26][26] ), .QN(n786) );
  SDFFNSRXL \regfile_reg[26][25]  ( .D(n3264), .SI(n788), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4472), .Q(\regfile[26][25] ), .QN(n787) );
  SDFFNSRXL \regfile_reg[26][24]  ( .D(n3262), .SI(n789), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4472), .Q(\regfile[26][24] ), .QN(n788) );
  SDFFNSRXL \regfile_reg[26][23]  ( .D(n3260), .SI(n790), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4472), .Q(\regfile[26][23] ), .QN(n789) );
  SDFFNSRXL \regfile_reg[26][22]  ( .D(n3258), .SI(n791), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4472), .Q(\regfile[26][22] ), .QN(n790) );
  SDFFNSRXL \regfile_reg[26][21]  ( .D(n3256), .SI(n792), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4472), .Q(\regfile[26][21] ), .QN(n791) );
  SDFFNSRXL \regfile_reg[26][20]  ( .D(n3254), .SI(n793), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4472), .Q(\regfile[26][20] ), .QN(n792) );
  SDFFNSRXL \regfile_reg[26][19]  ( .D(n3252), .SI(n794), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4472), .Q(\regfile[26][19] ), .QN(n793) );
  SDFFNSRXL \regfile_reg[26][18]  ( .D(n3250), .SI(n795), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4472), .Q(\regfile[26][18] ), .QN(n794) );
  SDFFNSRXL \regfile_reg[26][17]  ( .D(n3248), .SI(n796), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4472), .Q(\regfile[26][17] ), .QN(n795) );
  SDFFNSRXL \regfile_reg[26][16]  ( .D(n3246), .SI(n797), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4472), .Q(\regfile[26][16] ), .QN(n796) );
  SDFFNSRXL \regfile_reg[26][15]  ( .D(n3244), .SI(n798), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4472), .Q(\regfile[26][15] ), .QN(n797) );
  SDFFNSRXL \regfile_reg[26][14]  ( .D(n3242), .SI(n799), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4472), .Q(\regfile[26][14] ), .QN(n798) );
  SDFFNSRXL \regfile_reg[26][13]  ( .D(n3240), .SI(n800), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4472), .Q(\regfile[26][13] ), .QN(n799) );
  SDFFNSRXL \regfile_reg[26][12]  ( .D(n3238), .SI(n801), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4472), .Q(\regfile[26][12] ), .QN(n800) );
  SDFFNSRXL \regfile_reg[26][11]  ( .D(n3236), .SI(n802), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4472), .Q(\regfile[26][11] ), .QN(n801) );
  SDFFNSRXL \regfile_reg[26][10]  ( .D(n3234), .SI(n803), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4472), .Q(\regfile[26][10] ), .QN(n802) );
  SDFFNSRXL \regfile_reg[26][9]  ( .D(n3232), .SI(n804), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4473), .Q(\regfile[26][9] ), .QN(n803) );
  SDFFNSRXL \regfile_reg[26][8]  ( .D(n3230), .SI(n805), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4473), .Q(\regfile[26][8] ), .QN(n804) );
  SDFFNSRXL \regfile_reg[26][7]  ( .D(n3228), .SI(n806), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4473), .Q(\regfile[26][7] ), .QN(n805) );
  SDFFNSRXL \regfile_reg[26][6]  ( .D(n3226), .SI(n807), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4473), .Q(\regfile[26][6] ), .QN(n806) );
  SDFFNSRXL \regfile_reg[26][5]  ( .D(n3224), .SI(n808), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4473), .Q(\regfile[26][5] ), .QN(n807) );
  SDFFNSRXL \regfile_reg[26][4]  ( .D(n3222), .SI(n809), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4473), .Q(\regfile[26][4] ), .QN(n808) );
  SDFFNSRXL \regfile_reg[26][3]  ( .D(n3220), .SI(n810), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4473), .Q(\regfile[26][3] ), .QN(n809) );
  SDFFNSRXL \regfile_reg[26][2]  ( .D(n3218), .SI(n811), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4473), .Q(\regfile[26][2] ), .QN(n810) );
  SDFFNSRXL \regfile_reg[26][1]  ( .D(n3216), .SI(n812), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4473), .Q(\regfile[26][1] ), .QN(n811) );
  SDFFNSRXL \regfile_reg[26][0]  ( .D(n3214), .SI(n813), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4473), .Q(\regfile[26][0] ), .QN(n812) );
  SDFFNSRXL \regfile_reg[22][31]  ( .D(n3020), .SI(n910), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4478), .Q(\regfile[22][31] ), .QN(n909) );
  SDFFNSRXL \regfile_reg[22][30]  ( .D(n3018), .SI(n911), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4478), .Q(\regfile[22][30] ), .QN(n910) );
  SDFFNSRXL \regfile_reg[22][29]  ( .D(n3016), .SI(n912), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4479), .Q(\regfile[22][29] ), .QN(n911) );
  SDFFNSRXL \regfile_reg[22][28]  ( .D(n3014), .SI(n913), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4479), .Q(\regfile[22][28] ), .QN(n912) );
  SDFFNSRXL \regfile_reg[22][27]  ( .D(n3012), .SI(n914), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4479), .Q(\regfile[22][27] ), .QN(n913) );
  SDFFNSRXL \regfile_reg[22][26]  ( .D(n3010), .SI(n915), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4479), .Q(\regfile[22][26] ), .QN(n914) );
  SDFFNSRXL \regfile_reg[22][25]  ( .D(n3008), .SI(n916), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4479), .Q(\regfile[22][25] ), .QN(n915) );
  SDFFNSRXL \regfile_reg[22][24]  ( .D(n3006), .SI(n917), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4479), .Q(\regfile[22][24] ), .QN(n916) );
  SDFFNSRXL \regfile_reg[22][23]  ( .D(n3004), .SI(n918), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4479), .Q(\regfile[22][23] ), .QN(n917) );
  SDFFNSRXL \regfile_reg[22][22]  ( .D(n3002), .SI(n919), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4479), .Q(\regfile[22][22] ), .QN(n918) );
  SDFFNSRXL \regfile_reg[22][21]  ( .D(n3000), .SI(n920), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4479), .Q(\regfile[22][21] ), .QN(n919) );
  SDFFNSRXL \regfile_reg[22][20]  ( .D(n2998), .SI(n921), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4479), .Q(\regfile[22][20] ), .QN(n920) );
  SDFFNSRXL \regfile_reg[22][19]  ( .D(n2996), .SI(n922), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4479), .Q(\regfile[22][19] ), .QN(n921) );
  SDFFNSRXL \regfile_reg[22][18]  ( .D(n2994), .SI(n923), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4479), .Q(\regfile[22][18] ), .QN(n922) );
  SDFFNSRXL \regfile_reg[22][17]  ( .D(n2992), .SI(n924), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4479), .Q(\regfile[22][17] ), .QN(n923) );
  SDFFNSRXL \regfile_reg[22][16]  ( .D(n2990), .SI(n925), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4479), .Q(\regfile[22][16] ), .QN(n924) );
  SDFFNSRXL \regfile_reg[22][15]  ( .D(n2988), .SI(n926), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4479), .Q(\regfile[22][15] ), .QN(n925) );
  SDFFNSRXL \regfile_reg[22][14]  ( .D(n2986), .SI(n927), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4479), .Q(\regfile[22][14] ), .QN(n926) );
  SDFFNSRXL \regfile_reg[22][13]  ( .D(n2984), .SI(n928), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4479), .Q(\regfile[22][13] ), .QN(n927) );
  SDFFNSRXL \regfile_reg[22][12]  ( .D(n2982), .SI(n929), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4479), .Q(\regfile[22][12] ), .QN(n928) );
  SDFFNSRXL \regfile_reg[22][11]  ( .D(n2980), .SI(n930), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4480), .Q(\regfile[22][11] ), .QN(n929) );
  SDFFNSRXL \regfile_reg[22][10]  ( .D(n2978), .SI(n931), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4480), .Q(\regfile[22][10] ), .QN(n930) );
  SDFFNSRXL \regfile_reg[22][9]  ( .D(n2976), .SI(n932), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4480), .Q(\regfile[22][9] ), .QN(n931) );
  SDFFNSRXL \regfile_reg[22][8]  ( .D(n2974), .SI(n933), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4480), .Q(\regfile[22][8] ), .QN(n932) );
  SDFFNSRXL \regfile_reg[22][7]  ( .D(n2972), .SI(n934), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4480), .Q(\regfile[22][7] ), .QN(n933) );
  SDFFNSRXL \regfile_reg[22][6]  ( .D(n2970), .SI(n935), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4480), .Q(\regfile[22][6] ), .QN(n934) );
  SDFFNSRXL \regfile_reg[22][5]  ( .D(n2968), .SI(n936), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4480), .Q(\regfile[22][5] ), .QN(n935) );
  SDFFNSRXL \regfile_reg[22][4]  ( .D(n2966), .SI(n937), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4480), .Q(\regfile[22][4] ), .QN(n936) );
  SDFFNSRXL \regfile_reg[22][3]  ( .D(n2964), .SI(n938), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4480), .Q(\regfile[22][3] ), .QN(n937) );
  SDFFNSRXL \regfile_reg[22][2]  ( .D(n2962), .SI(n939), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4480), .Q(\regfile[22][2] ), .QN(n938) );
  SDFFNSRXL \regfile_reg[22][1]  ( .D(n2960), .SI(n940), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4480), .Q(\regfile[22][1] ), .QN(n939) );
  SDFFNSRXL \regfile_reg[22][0]  ( .D(n2958), .SI(n941), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4480), .Q(\regfile[22][0] ), .QN(n940) );
  SDFFNSRXL \regfile_reg[18][31]  ( .D(n2764), .SI(n1038), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4486), .Q(\regfile[18][31] ), .QN(n1037) );
  SDFFNSRXL \regfile_reg[18][30]  ( .D(n2762), .SI(n1039), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4486), .Q(\regfile[18][30] ), .QN(n1038) );
  SDFFNSRXL \regfile_reg[18][29]  ( .D(n2760), .SI(n1040), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4486), .Q(\regfile[18][29] ), .QN(n1039) );
  SDFFNSRXL \regfile_reg[18][28]  ( .D(n2758), .SI(n1041), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4486), .Q(\regfile[18][28] ), .QN(n1040) );
  SDFFNSRXL \regfile_reg[18][27]  ( .D(n2756), .SI(n1042), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4486), .Q(\regfile[18][27] ), .QN(n1041) );
  SDFFNSRXL \regfile_reg[18][26]  ( .D(n2754), .SI(n1043), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4486), .Q(\regfile[18][26] ), .QN(n1042) );
  SDFFNSRXL \regfile_reg[18][25]  ( .D(n2752), .SI(n1044), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4486), .Q(\regfile[18][25] ), .QN(n1043) );
  SDFFNSRXL \regfile_reg[18][24]  ( .D(n2750), .SI(n1045), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4486), .Q(\regfile[18][24] ), .QN(n1044) );
  SDFFNSRXL \regfile_reg[18][23]  ( .D(n2748), .SI(n1046), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4486), .Q(\regfile[18][23] ), .QN(n1045) );
  SDFFNSRXL \regfile_reg[18][22]  ( .D(n2746), .SI(n1047), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4486), .Q(\regfile[18][22] ), .QN(n1046) );
  SDFFNSRXL \regfile_reg[18][21]  ( .D(n2744), .SI(n1048), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4486), .Q(\regfile[18][21] ), .QN(n1047) );
  SDFFNSRXL \regfile_reg[18][20]  ( .D(n2742), .SI(n1049), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4486), .Q(\regfile[18][20] ), .QN(n1048) );
  SDFFNSRXL \regfile_reg[18][19]  ( .D(n2740), .SI(n1050), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4486), .Q(\regfile[18][19] ), .QN(n1049) );
  SDFFNSRXL \regfile_reg[18][18]  ( .D(n2738), .SI(n1051), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4486), .Q(\regfile[18][18] ), .QN(n1050) );
  SDFFNSRXL \regfile_reg[18][17]  ( .D(n2736), .SI(n1052), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4486), .Q(\regfile[18][17] ), .QN(n1051) );
  SDFFNSRXL \regfile_reg[18][16]  ( .D(n2734), .SI(n1053), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4486), .Q(\regfile[18][16] ), .QN(n1052) );
  SDFFNSRXL \regfile_reg[18][15]  ( .D(n2732), .SI(n1054), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4486), .Q(\regfile[18][15] ), .QN(n1053) );
  SDFFNSRXL \regfile_reg[18][14]  ( .D(n2730), .SI(n1055), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4486), .Q(\regfile[18][14] ), .QN(n1054) );
  SDFFNSRXL \regfile_reg[18][13]  ( .D(n2728), .SI(n1056), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4487), .Q(\regfile[18][13] ), .QN(n1055) );
  SDFFNSRXL \regfile_reg[18][12]  ( .D(n2726), .SI(n1057), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4487), .Q(\regfile[18][12] ), .QN(n1056) );
  SDFFNSRXL \regfile_reg[18][11]  ( .D(n2724), .SI(n1058), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4487), .Q(\regfile[18][11] ), .QN(n1057) );
  SDFFNSRXL \regfile_reg[18][10]  ( .D(n2722), .SI(n1059), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4487), .Q(\regfile[18][10] ), .QN(n1058) );
  SDFFNSRXL \regfile_reg[18][9]  ( .D(n2720), .SI(n1060), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4487), .Q(\regfile[18][9] ), .QN(n1059) );
  SDFFNSRXL \regfile_reg[18][8]  ( .D(n2718), .SI(n1061), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4487), .Q(\regfile[18][8] ), .QN(n1060) );
  SDFFNSRXL \regfile_reg[18][7]  ( .D(n2716), .SI(n1062), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4487), .Q(\regfile[18][7] ), .QN(n1061) );
  SDFFNSRXL \regfile_reg[18][6]  ( .D(n2714), .SI(n1063), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4487), .Q(\regfile[18][6] ), .QN(n1062) );
  SDFFNSRXL \regfile_reg[18][5]  ( .D(n2712), .SI(n1064), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4487), .Q(\regfile[18][5] ), .QN(n1063) );
  SDFFNSRXL \regfile_reg[18][4]  ( .D(n2710), .SI(n1065), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4487), .Q(\regfile[18][4] ), .QN(n1064) );
  SDFFNSRXL \regfile_reg[18][3]  ( .D(n2708), .SI(n1066), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4487), .Q(\regfile[18][3] ), .QN(n1065) );
  SDFFNSRXL \regfile_reg[18][2]  ( .D(n2706), .SI(n1067), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4487), .Q(\regfile[18][2] ), .QN(n1066) );
  SDFFNSRXL \regfile_reg[18][1]  ( .D(n2704), .SI(n1068), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4487), .Q(\regfile[18][1] ), .QN(n1067) );
  SDFFNSRXL \regfile_reg[18][0]  ( .D(n2702), .SI(n1069), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4487), .Q(\regfile[18][0] ), .QN(n1068) );
  SDFFNSRXL \regfile_reg[14][31]  ( .D(n2508), .SI(n1166), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4493), .Q(\regfile[14][31] ), .QN(n1165) );
  SDFFNSRXL \regfile_reg[14][30]  ( .D(n2506), .SI(n1167), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4493), .Q(\regfile[14][30] ), .QN(n1166) );
  SDFFNSRXL \regfile_reg[14][29]  ( .D(n2504), .SI(n1168), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4493), .Q(\regfile[14][29] ), .QN(n1167) );
  SDFFNSRXL \regfile_reg[14][28]  ( .D(n2502), .SI(n1169), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4493), .Q(\regfile[14][28] ), .QN(n1168) );
  SDFFNSRXL \regfile_reg[14][27]  ( .D(n2500), .SI(n1170), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4493), .Q(\regfile[14][27] ), .QN(n1169) );
  SDFFNSRXL \regfile_reg[14][26]  ( .D(n2498), .SI(n1171), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4493), .Q(\regfile[14][26] ), .QN(n1170) );
  SDFFNSRXL \regfile_reg[14][25]  ( .D(n2496), .SI(n1172), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4493), .Q(\regfile[14][25] ), .QN(n1171) );
  SDFFNSRXL \regfile_reg[14][24]  ( .D(n2494), .SI(n1173), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4493), .Q(\regfile[14][24] ), .QN(n1172) );
  SDFFNSRXL \regfile_reg[14][23]  ( .D(n2492), .SI(n1174), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4493), .Q(\regfile[14][23] ), .QN(n1173) );
  SDFFNSRXL \regfile_reg[14][22]  ( .D(n2490), .SI(n1175), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4493), .Q(\regfile[14][22] ), .QN(n1174) );
  SDFFNSRXL \regfile_reg[14][21]  ( .D(n2488), .SI(n1176), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4493), .Q(\regfile[14][21] ), .QN(n1175) );
  SDFFNSRXL \regfile_reg[14][20]  ( .D(n2486), .SI(n1177), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4493), .Q(\regfile[14][20] ), .QN(n1176) );
  SDFFNSRXL \regfile_reg[14][19]  ( .D(n2484), .SI(n1178), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4493), .Q(\regfile[14][19] ), .QN(n1177) );
  SDFFNSRXL \regfile_reg[14][18]  ( .D(n2482), .SI(n1179), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4493), .Q(\regfile[14][18] ), .QN(n1178) );
  SDFFNSRXL \regfile_reg[14][17]  ( .D(n2480), .SI(n1180), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4493), .Q(\regfile[14][17] ), .QN(n1179) );
  SDFFNSRXL \regfile_reg[14][16]  ( .D(n2478), .SI(n1181), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4493), .Q(\regfile[14][16] ), .QN(n1180) );
  SDFFNSRXL \regfile_reg[14][15]  ( .D(n2476), .SI(n1182), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4494), .Q(\regfile[14][15] ), .QN(n1181) );
  SDFFNSRXL \regfile_reg[14][14]  ( .D(n2474), .SI(n1183), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4494), .Q(\regfile[14][14] ), .QN(n1182) );
  SDFFNSRXL \regfile_reg[14][13]  ( .D(n2472), .SI(n1184), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4494), .Q(\regfile[14][13] ), .QN(n1183) );
  SDFFNSRXL \regfile_reg[14][12]  ( .D(n2470), .SI(n1185), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4494), .Q(\regfile[14][12] ), .QN(n1184) );
  SDFFNSRXL \regfile_reg[14][11]  ( .D(n2468), .SI(n1186), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4494), .Q(\regfile[14][11] ), .QN(n1185) );
  SDFFNSRXL \regfile_reg[14][10]  ( .D(n2466), .SI(n1187), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4494), .Q(\regfile[14][10] ), .QN(n1186) );
  SDFFNSRXL \regfile_reg[14][9]  ( .D(n2464), .SI(n1188), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4494), .Q(\regfile[14][9] ), .QN(n1187) );
  SDFFNSRXL \regfile_reg[14][8]  ( .D(n2462), .SI(n1189), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4494), .Q(\regfile[14][8] ), .QN(n1188) );
  SDFFNSRXL \regfile_reg[14][7]  ( .D(n2460), .SI(n1190), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4494), .Q(\regfile[14][7] ), .QN(n1189) );
  SDFFNSRXL \regfile_reg[14][6]  ( .D(n2458), .SI(n1191), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4494), .Q(\regfile[14][6] ), .QN(n1190) );
  SDFFNSRXL \regfile_reg[14][5]  ( .D(n2456), .SI(n1192), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4494), .Q(\regfile[14][5] ), .QN(n1191) );
  SDFFNSRXL \regfile_reg[14][4]  ( .D(n2454), .SI(n1193), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4494), .Q(\regfile[14][4] ), .QN(n1192) );
  SDFFNSRXL \regfile_reg[14][3]  ( .D(n2452), .SI(n1194), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4494), .Q(\regfile[14][3] ), .QN(n1193) );
  SDFFNSRXL \regfile_reg[14][2]  ( .D(n2450), .SI(n1195), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4494), .Q(\regfile[14][2] ), .QN(n1194) );
  SDFFNSRXL \regfile_reg[14][1]  ( .D(n2448), .SI(n1196), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4494), .Q(\regfile[14][1] ), .QN(n1195) );
  SDFFNSRXL \regfile_reg[14][0]  ( .D(n2446), .SI(n1197), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4494), .Q(\regfile[14][0] ), .QN(n1196) );
  SDFFNSRXL \regfile_reg[10][31]  ( .D(n2252), .SI(n1294), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4500), .Q(\regfile[10][31] ), .QN(n1293) );
  SDFFNSRXL \regfile_reg[10][30]  ( .D(n2250), .SI(n1295), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4500), .Q(\regfile[10][30] ), .QN(n1294) );
  SDFFNSRXL \regfile_reg[10][29]  ( .D(n2248), .SI(n1296), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4500), .Q(\regfile[10][29] ), .QN(n1295) );
  SDFFNSRXL \regfile_reg[10][28]  ( .D(n2246), .SI(n1297), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4500), .Q(\regfile[10][28] ), .QN(n1296) );
  SDFFNSRXL \regfile_reg[10][27]  ( .D(n2244), .SI(n1298), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4500), .Q(\regfile[10][27] ), .QN(n1297) );
  SDFFNSRXL \regfile_reg[10][26]  ( .D(n2242), .SI(n1299), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4500), .Q(\regfile[10][26] ), .QN(n1298) );
  SDFFNSRXL \regfile_reg[10][25]  ( .D(n2240), .SI(n1300), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4500), .Q(\regfile[10][25] ), .QN(n1299) );
  SDFFNSRXL \regfile_reg[10][24]  ( .D(n2238), .SI(n1301), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4500), .Q(\regfile[10][24] ), .QN(n1300) );
  SDFFNSRXL \regfile_reg[10][23]  ( .D(n2236), .SI(n1302), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4500), .Q(\regfile[10][23] ), .QN(n1301) );
  SDFFNSRXL \regfile_reg[10][22]  ( .D(n2234), .SI(n1303), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4500), .Q(\regfile[10][22] ), .QN(n1302) );
  SDFFNSRXL \regfile_reg[10][21]  ( .D(n2232), .SI(n1304), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4500), .Q(\regfile[10][21] ), .QN(n1303) );
  SDFFNSRXL \regfile_reg[10][20]  ( .D(n2230), .SI(n1305), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4500), .Q(\regfile[10][20] ), .QN(n1304) );
  SDFFNSRXL \regfile_reg[10][19]  ( .D(n2228), .SI(n1306), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4500), .Q(\regfile[10][19] ), .QN(n1305) );
  SDFFNSRXL \regfile_reg[10][18]  ( .D(n2226), .SI(n1307), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4500), .Q(\regfile[10][18] ), .QN(n1306) );
  SDFFNSRXL \regfile_reg[10][17]  ( .D(n2224), .SI(n1308), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4501), .Q(\regfile[10][17] ), .QN(n1307) );
  SDFFNSRXL \regfile_reg[10][16]  ( .D(n2222), .SI(n1309), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4501), .Q(\regfile[10][16] ), .QN(n1308) );
  SDFFNSRXL \regfile_reg[10][15]  ( .D(n2220), .SI(n1310), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4501), .Q(\regfile[10][15] ), .QN(n1309) );
  SDFFNSRXL \regfile_reg[10][14]  ( .D(n2218), .SI(n1311), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4501), .Q(\regfile[10][14] ), .QN(n1310) );
  SDFFNSRXL \regfile_reg[10][13]  ( .D(n2216), .SI(n1312), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4501), .Q(\regfile[10][13] ), .QN(n1311) );
  SDFFNSRXL \regfile_reg[10][12]  ( .D(n2214), .SI(n1313), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4501), .Q(\regfile[10][12] ), .QN(n1312) );
  SDFFNSRXL \regfile_reg[10][11]  ( .D(n2212), .SI(n1314), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4501), .Q(\regfile[10][11] ), .QN(n1313) );
  SDFFNSRXL \regfile_reg[10][10]  ( .D(n2210), .SI(n1315), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4501), .Q(\regfile[10][10] ), .QN(n1314) );
  SDFFNSRXL \regfile_reg[10][9]  ( .D(n2208), .SI(n1316), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4501), .Q(\regfile[10][9] ), .QN(n1315) );
  SDFFNSRXL \regfile_reg[10][8]  ( .D(n2206), .SI(n1317), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4501), .Q(\regfile[10][8] ), .QN(n1316) );
  SDFFNSRXL \regfile_reg[10][7]  ( .D(n2204), .SI(n1318), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4501), .Q(\regfile[10][7] ), .QN(n1317) );
  SDFFNSRXL \regfile_reg[10][6]  ( .D(n2202), .SI(n1319), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4501), .Q(\regfile[10][6] ), .QN(n1318) );
  SDFFNSRXL \regfile_reg[10][5]  ( .D(n2200), .SI(n1320), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4501), .Q(\regfile[10][5] ), .QN(n1319) );
  SDFFNSRXL \regfile_reg[10][4]  ( .D(n2198), .SI(n1321), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4501), .Q(\regfile[10][4] ), .QN(n1320) );
  SDFFNSRXL \regfile_reg[10][3]  ( .D(n2196), .SI(n1322), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4501), .Q(\regfile[10][3] ), .QN(n1321) );
  SDFFNSRXL \regfile_reg[10][2]  ( .D(n2194), .SI(n1323), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4501), .Q(\regfile[10][2] ), .QN(n1322) );
  SDFFNSRXL \regfile_reg[10][1]  ( .D(n2192), .SI(n1324), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4501), .Q(\regfile[10][1] ), .QN(n1323) );
  SDFFNSRXL \regfile_reg[10][0]  ( .D(n2190), .SI(n1325), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4501), .Q(\regfile[10][0] ), .QN(n1324) );
  SDFFNSRXL \regfile_reg[6][31]  ( .D(n1996), .SI(n1422), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4507), .Q(\regfile[6][31] ), .QN(n1421) );
  SDFFNSRXL \regfile_reg[6][30]  ( .D(n1994), .SI(n1423), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4507), .Q(\regfile[6][30] ), .QN(n1422) );
  SDFFNSRXL \regfile_reg[6][29]  ( .D(n1992), .SI(n1424), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4507), .Q(\regfile[6][29] ), .QN(n1423) );
  SDFFNSRXL \regfile_reg[6][28]  ( .D(n1990), .SI(n1425), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4507), .Q(\regfile[6][28] ), .QN(n1424) );
  SDFFNSRXL \regfile_reg[6][27]  ( .D(n1988), .SI(n1426), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4507), .Q(\regfile[6][27] ), .QN(n1425) );
  SDFFNSRXL \regfile_reg[6][26]  ( .D(n1986), .SI(n1427), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4507), .Q(\regfile[6][26] ), .QN(n1426) );
  SDFFNSRXL \regfile_reg[6][25]  ( .D(n1984), .SI(n1428), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4507), .Q(\regfile[6][25] ), .QN(n1427) );
  SDFFNSRXL \regfile_reg[6][24]  ( .D(n1982), .SI(n1429), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4507), .Q(\regfile[6][24] ), .QN(n1428) );
  SDFFNSRXL \regfile_reg[6][23]  ( .D(n1980), .SI(n1430), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4507), .Q(\regfile[6][23] ), .QN(n1429) );
  SDFFNSRXL \regfile_reg[6][22]  ( .D(n1978), .SI(n1431), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4507), .Q(\regfile[6][22] ), .QN(n1430) );
  SDFFNSRXL \regfile_reg[6][21]  ( .D(n1976), .SI(n1432), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4507), .Q(\regfile[6][21] ), .QN(n1431) );
  SDFFNSRXL \regfile_reg[6][20]  ( .D(n1974), .SI(n1433), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4507), .Q(\regfile[6][20] ), .QN(n1432) );
  SDFFNSRXL \regfile_reg[6][19]  ( .D(n1972), .SI(n1434), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4508), .Q(\regfile[6][19] ), .QN(n1433) );
  SDFFNSRXL \regfile_reg[6][18]  ( .D(n1970), .SI(n1435), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4508), .Q(\regfile[6][18] ), .QN(n1434) );
  SDFFNSRXL \regfile_reg[6][17]  ( .D(n1968), .SI(n1436), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4508), .Q(\regfile[6][17] ), .QN(n1435) );
  SDFFNSRXL \regfile_reg[6][16]  ( .D(n1966), .SI(n1437), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4508), .Q(\regfile[6][16] ), .QN(n1436) );
  SDFFNSRXL \regfile_reg[6][15]  ( .D(n1964), .SI(n1438), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4508), .Q(\regfile[6][15] ), .QN(n1437) );
  SDFFNSRXL \regfile_reg[6][14]  ( .D(n1962), .SI(n1439), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4508), .Q(\regfile[6][14] ), .QN(n1438) );
  SDFFNSRXL \regfile_reg[6][13]  ( .D(n1960), .SI(n1440), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4508), .Q(\regfile[6][13] ), .QN(n1439) );
  SDFFNSRXL \regfile_reg[6][12]  ( .D(n1958), .SI(n1441), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4508), .Q(\regfile[6][12] ), .QN(n1440) );
  SDFFNSRXL \regfile_reg[6][11]  ( .D(n1956), .SI(n1442), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4508), .Q(\regfile[6][11] ), .QN(n1441) );
  SDFFNSRXL \regfile_reg[6][10]  ( .D(n1954), .SI(n1443), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4508), .Q(\regfile[6][10] ), .QN(n1442) );
  SDFFNSRXL \regfile_reg[6][9]  ( .D(n1952), .SI(n1444), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4508), .Q(\regfile[6][9] ), .QN(n1443) );
  SDFFNSRXL \regfile_reg[6][8]  ( .D(n1950), .SI(n1445), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4508), .Q(\regfile[6][8] ), .QN(n1444) );
  SDFFNSRXL \regfile_reg[6][7]  ( .D(n1948), .SI(n1446), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4508), .Q(\regfile[6][7] ), .QN(n1445) );
  SDFFNSRXL \regfile_reg[6][6]  ( .D(n1946), .SI(n1447), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4508), .Q(\regfile[6][6] ), .QN(n1446) );
  SDFFNSRXL \regfile_reg[6][5]  ( .D(n1944), .SI(n1448), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4508), .Q(\regfile[6][5] ), .QN(n1447) );
  SDFFNSRXL \regfile_reg[6][4]  ( .D(n1942), .SI(n1449), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4508), .Q(\regfile[6][4] ), .QN(n1448) );
  SDFFNSRXL \regfile_reg[6][3]  ( .D(n1940), .SI(n1450), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4508), .Q(\regfile[6][3] ), .QN(n1449) );
  SDFFNSRXL \regfile_reg[6][2]  ( .D(n1938), .SI(n1451), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4508), .Q(\regfile[6][2] ), .QN(n1450) );
  SDFFNSRXL \regfile_reg[6][1]  ( .D(n1936), .SI(n1452), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4509), .Q(\regfile[6][1] ), .QN(n1451) );
  SDFFNSRXL \regfile_reg[6][0]  ( .D(n1934), .SI(n1453), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4509), .Q(\regfile[6][0] ), .QN(n1452) );
  SDFFNSRXL \regfile_reg[3][31]  ( .D(n1804), .SI(n1518), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4512), .Q(\regfile[3][31] ), .QN(n1517) );
  SDFFNSRXL \regfile_reg[3][30]  ( .D(n1802), .SI(n1519), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4512), .Q(\regfile[3][30] ), .QN(n1518) );
  SDFFNSRXL \regfile_reg[3][29]  ( .D(n1800), .SI(n1520), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4512), .Q(\regfile[3][29] ), .QN(n1519) );
  SDFFNSRXL \regfile_reg[3][28]  ( .D(n1798), .SI(n1521), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4512), .Q(\regfile[3][28] ), .QN(n1520) );
  SDFFNSRXL \regfile_reg[3][27]  ( .D(n1796), .SI(n1522), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4512), .Q(\regfile[3][27] ), .QN(n1521) );
  SDFFNSRXL \regfile_reg[3][26]  ( .D(n1794), .SI(n1523), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4512), .Q(\regfile[3][26] ), .QN(n1522) );
  SDFFNSRXL \regfile_reg[3][25]  ( .D(n1792), .SI(n1524), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4513), .Q(\regfile[3][25] ), .QN(n1523) );
  SDFFNSRXL \regfile_reg[3][24]  ( .D(n1790), .SI(n1525), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4513), .Q(\regfile[3][24] ), .QN(n1524) );
  SDFFNSRXL \regfile_reg[3][22]  ( .D(n1786), .SI(n1527), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4513), .Q(\regfile[3][22] ), .QN(n1526) );
  SDFFNSRXL \regfile_reg[3][21]  ( .D(n1784), .SI(n1528), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4513), .Q(\regfile[3][21] ), .QN(n1527) );
  SDFFNSRXL \regfile_reg[3][15]  ( .D(n1772), .SI(n1534), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4513), .Q(\regfile[3][15] ), .QN(n1533) );
  SDFFNSRXL \regfile_reg[3][14]  ( .D(n1770), .SI(n1535), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4513), .Q(\regfile[3][14] ), .QN(n1534) );
  SDFFNSRXL \regfile_reg[3][13]  ( .D(n1768), .SI(n1536), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4513), .Q(\regfile[3][13] ), .QN(n1535) );
  SDFFNSRXL \regfile_reg[3][12]  ( .D(n1766), .SI(n1537), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4513), .Q(\regfile[3][12] ), .QN(n1536) );
  SDFFNSRXL \regfile_reg[3][11]  ( .D(n1764), .SI(n1895), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4513), .Q(\regfile[3][11] ), .QN(n1537) );
  SDFFNSRXL \regfile_reg[3][9]  ( .D(n1760), .SI(n1540), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4513), .Q(\regfile[3][9] ), .QN(n1539) );
  SDFFNSRXL \regfile_reg[3][8]  ( .D(n1758), .SI(n1541), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4513), .Q(\regfile[3][8] ), .QN(n1540) );
  SDFFNSRXL \regfile_reg[3][5]  ( .D(n1752), .SI(n1544), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4514), .Q(\regfile[3][5] ), .QN(n1543) );
  SDFFNSRXL \regfile_reg[3][1]  ( .D(n1744), .SI(n1548), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4514), .Q(\regfile[3][1] ), .QN(n1547) );
  SDFFNSRXL \regfile_reg[1][31]  ( .D(n1676), .SI(n1783), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4516), .Q(\regfile[1][31] ), .QN(n1581) );
  SDFFNSRXL \regfile_reg[1][30]  ( .D(n1674), .SI(n1583), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4516), .Q(\regfile[1][30] ), .QN(n1582) );
  SDFFNSRXL \regfile_reg[1][29]  ( .D(n1672), .SI(n1584), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4516), .Q(\regfile[1][29] ), .QN(n1583) );
  SDFFNSRXL \regfile_reg[1][28]  ( .D(n1670), .SI(n1585), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4516), .Q(\regfile[1][28] ), .QN(n1584) );
  SDFFNSRXL \regfile_reg[1][27]  ( .D(n1668), .SI(n1586), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4516), .Q(\regfile[1][27] ), .QN(n1585) );
  SDFFNSRXL \regfile_reg[1][26]  ( .D(n1666), .SI(n1587), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4516), .Q(\regfile[1][26] ), .QN(n1586) );
  SDFFNSRXL \regfile_reg[1][25]  ( .D(n1664), .SI(n1767), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4516), .Q(\regfile[1][25] ), .QN(n1587) );
  SDFFNSRXL \regfile_reg[1][24]  ( .D(n1662), .SI(n1589), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4516), .Q(\regfile[1][24] ), .QN(n1588) );
  SDFFNSRXL \regfile_reg[1][23]  ( .D(n1660), .SI(n1590), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4516), .Q(\regfile[1][23] ), .QN(n1589) );
  SDFFNSRXL \regfile_reg[1][22]  ( .D(n1658), .SI(n1591), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4516), .Q(\regfile[1][22] ), .QN(n1590) );
  SDFFNSRXL \regfile_reg[1][21]  ( .D(n1656), .SI(n1592), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4516), .Q(\regfile[1][21] ), .QN(n1591) );
  SDFFNSRXL \regfile_reg[1][20]  ( .D(n1654), .SI(n1775), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4516), .Q(\regfile[1][20] ), .QN(n1592) );
  SDFFNSRXL \regfile_reg[1][19]  ( .D(n1652), .SI(n1594), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4516), .Q(\regfile[1][19] ), .QN(n1593) );
  SDFFNSRXL \regfile_reg[1][18]  ( .D(n1650), .SI(n1595), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4516), .Q(\regfile[1][18] ), .QN(n1594) );
  SDFFNSRXL \regfile_reg[1][17]  ( .D(n1648), .SI(n1596), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4517), .Q(\regfile[1][17] ), .QN(n1595) );
  SDFFNSRXL \regfile_reg[1][16]  ( .D(n1646), .SI(n1597), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4517), .Q(\regfile[1][16] ), .QN(n1596) );
  SDFFNSRXL \regfile_reg[1][15]  ( .D(n1644), .SI(n1598), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4517), .Q(\regfile[1][15] ), .QN(n1597) );
  SDFFNSRXL \regfile_reg[1][14]  ( .D(n1642), .SI(n1599), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4517), .Q(\regfile[1][14] ), .QN(n1598) );
  SDFFNSRXL \regfile_reg[1][13]  ( .D(n1640), .SI(n1600), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4517), .Q(\regfile[1][13] ), .QN(n1599) );
  SDFFNSRXL \regfile_reg[1][12]  ( .D(n1638), .SI(n1601), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4517), .Q(\regfile[1][12] ), .QN(n1600) );
  SDFFNSRXL \regfile_reg[1][11]  ( .D(n1636), .SI(n1602), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4517), .Q(\regfile[1][11] ), .QN(n1601) );
  SDFFNSRXL \regfile_reg[1][10]  ( .D(n1634), .SI(n1773), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4517), .Q(\regfile[1][10] ), .QN(n1602) );
  SDFFNSRXL \regfile_reg[1][9]  ( .D(n1632), .SI(n1765), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4517), .Q(\regfile[1][9] ), .QN(n1603) );
  SDFFNSRXL \regfile_reg[1][8]  ( .D(n1630), .SI(n1605), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4517), .Q(\regfile[1][8] ), .QN(n1604) );
  SDFFNSRXL \regfile_reg[1][7]  ( .D(n1628), .SI(n1606), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4517), .Q(\regfile[1][7] ), .QN(n1605) );
  SDFFNSRXL \regfile_reg[1][6]  ( .D(n1626), .SI(n1763), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4517), .Q(\regfile[1][6] ), .QN(n1606) );
  SDFFNSRXL \regfile_reg[1][5]  ( .D(n1624), .SI(n1771), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4517), .Q(\regfile[1][5] ), .QN(n1607) );
  SDFFNSRXL \regfile_reg[1][4]  ( .D(n1622), .SI(n1769), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4517), .Q(\regfile[1][4] ), .QN(n1608) );
  SDFFNSRXL \regfile_reg[1][3]  ( .D(n1620), .SI(n1759), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4517), .Q(\regfile[1][3] ), .QN(n1609) );
  SDFFNSRXL \regfile_reg[1][2]  ( .D(n1618), .SI(n1611), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4517), .Q(\regfile[1][2] ), .QN(n1610) );
  SDFFNSRXL \regfile_reg[1][1]  ( .D(n1616), .SI(n1757), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4517), .Q(\regfile[1][1] ), .QN(n1611) );
  SDFFNSRXL \regfile_reg[1][0]  ( .D(n1614), .SI(test_si1), .SE(test_se), 
        .CKN(clk), .SN(1'b1), .RN(n4517), .Q(\regfile[1][0] ), .QN(n1612) );
  SDFFRXL \EX_reg[2]  ( .D(n3607), .SI(n638), .SE(test_se), .CK(clk), .RN(
        n4451), .Q(n1943), .QN(n639) );
  SDFFRXL \Immediate_SE_reg[1]  ( .D(n142), .SI(n601), .SE(test_se), .CK(clk), 
        .RN(n4462), .Q(n1951), .QN(n612) );
  SDFFRXL \RData2_reg[16]  ( .D(next_RData2[16]), .SI(n1655), .SE(test_se), 
        .CK(clk), .RN(n4458), .Q(RData2[16]), .QN(n1667) );
  SDFFRXL \RData2_reg[4]  ( .D(next_RData2[4]), .SI(n1647), .SE(test_se), .CK(
        clk), .RN(n4459), .Q(RData2[4]), .QN(n1665) );
  SDFFRXL \RData2_reg[14]  ( .D(next_RData2[14]), .SI(n1641), .SE(test_se), 
        .CK(clk), .RN(n4458), .Q(RData2[14]), .QN(n1663) );
  SDFFRXL \RData2_reg[0]  ( .D(next_RData2[0]), .SI(n1617), .SE(test_se), .CK(
        clk), .RN(n4459), .Q(RData2[0]), .QN(n1661) );
  SDFFRXL \RData2_reg[12]  ( .D(next_RData2[12]), .SI(n1619), .SE(test_se), 
        .CK(clk), .RN(n4458), .Q(RData2[12]), .QN(n1659) );
  SDFFRXL \RData2_reg[1]  ( .D(next_RData2[1]), .SI(n1661), .SE(test_se), .CK(
        clk), .RN(n4459), .Q(RData2[1]), .QN(n1657) );
  SDFFRXL \RData2_reg[15]  ( .D(next_RData2[15]), .SI(n1663), .SE(test_se), 
        .CK(clk), .RN(n4458), .Q(RData2[15]), .QN(n1655) );
  SDFFRXL \RData2_reg[5]  ( .D(next_RData2[5]), .SI(n1665), .SE(test_se), .CK(
        clk), .RN(n4459), .Q(RData2[5]), .QN(n1653) );
  SDFFRXL \RData2_reg[7]  ( .D(next_RData2[7]), .SI(n1649), .SE(test_se), .CK(
        clk), .RN(n4459), .Q(RData2[7]), .QN(n1651) );
  SDFFRXL \RData2_reg[6]  ( .D(next_RData2[6]), .SI(n1653), .SE(test_se), .CK(
        clk), .RN(n4459), .Q(RData2[6]), .QN(n1649) );
  SDFFRXL \RData2_reg[3]  ( .D(next_RData2[3]), .SI(n1645), .SE(test_se), .CK(
        clk), .RN(n4459), .Q(RData2[3]), .QN(n1647) );
  SDFFRXL \RData2_reg[2]  ( .D(next_RData2[2]), .SI(n1657), .SE(test_se), .CK(
        clk), .RN(n4459), .Q(RData2[2]), .QN(n1645) );
  SDFFRXL \RData2_reg[10]  ( .D(next_RData2[10]), .SI(n1637), .SE(test_se), 
        .CK(clk), .RN(n4458), .Q(RData2[10]), .QN(n1643) );
  SDFFRXL \RData2_reg[13]  ( .D(next_RData2[13]), .SI(n1659), .SE(test_se), 
        .CK(clk), .RN(n4458), .Q(RData2[13]), .QN(n1641) );
  SDFFRXL \RData2_reg[8]  ( .D(next_RData2[8]), .SI(n1651), .SE(test_se), .CK(
        clk), .RN(n4459), .Q(RData2[8]), .QN(n1639) );
  SDFFRXL \RData2_reg[9]  ( .D(next_RData2[9]), .SI(n1639), .SE(test_se), .CK(
        clk), .RN(n4459), .Q(RData2[9]), .QN(n1637) );
  SDFFRXL \RData1_reg[0]  ( .D(next_RData1[0]), .SI(n1901), .SE(test_se), .CK(
        clk), .RN(n4457), .Q(RData1[0]), .QN(n1635) );
  SDFFRXL \RData1_reg[8]  ( .D(next_RData1[8]), .SI(n44), .SE(test_se), .CK(
        clk), .RN(n4456), .Q(RData1[8]), .QN(n1633) );
  SDFFRXL \RData1_reg[4]  ( .D(next_RData1[4]), .SI(n41), .SE(test_se), .CK(
        clk), .RN(n4456), .Q(RData1[4]), .QN(n1631) );
  SDFFRXL \RData1_reg[10]  ( .D(next_RData1[10]), .SI(n45), .SE(test_se), .CK(
        clk), .RN(n4456), .Q(RData1[10]), .QN(n1629) );
  SDFFRXL \RData1_reg[12]  ( .D(next_RData1[12]), .SI(n46), .SE(test_se), .CK(
        clk), .RN(n4456), .Q(RData1[12]), .QN(n1627) );
  SDFFRXL \RData1_reg[14]  ( .D(next_RData1[14]), .SI(n70), .SE(test_se), .CK(
        clk), .RN(n4455), .Q(RData1[14]), .QN(n1625) );
  SDFFRXL \RData2_reg[25]  ( .D(next_RData2[25]), .SI(n1621), .SE(test_se), 
        .CK(clk), .RN(n4457), .Q(RData2[25]), .QN(n1623) );
  SDFFRXL \RData2_reg[24]  ( .D(next_RData2[24]), .SI(n59), .SE(test_se), .CK(
        clk), .RN(n4457), .Q(RData2[24]), .QN(n1621) );
  SDFFRXL \RData2_reg[11]  ( .D(next_RData2[11]), .SI(n1643), .SE(test_se), 
        .CK(clk), .RN(n4458), .Q(RData2[11]), .QN(n1619) );
  SDFFRXL \RData1_reg[31]  ( .D(next_RData1[31]), .SI(n1615), .SE(test_se), 
        .CK(clk), .RN(n4454), .Q(RData1[31]), .QN(n1617) );
  SDFFRXL \RData1_reg[30]  ( .D(next_RData1[30]), .SI(n1613), .SE(test_se), 
        .CK(clk), .RN(n4454), .Q(RData1[30]), .QN(n1615) );
  SDFFRXL \RData1_reg[29]  ( .D(next_RData1[29]), .SI(n101), .SE(test_se), 
        .CK(clk), .RN(n4454), .Q(RData1[29]), .QN(n1613) );
  SDFFRXL \RData1_reg[28]  ( .D(next_RData1[28]), .SI(n84), .SE(test_se), .CK(
        clk), .RN(n4454), .Q(RData1[28]), .QN(n101) );
  SDFFRXL \RData1_reg[27]  ( .D(next_RData1[27]), .SI(n80), .SE(test_se), .CK(
        clk), .RN(n4454), .Q(RData1[27]), .QN(n84) );
  SDFFRXL \RData2_reg[29]  ( .D(next_RData2[29]), .SI(n81), .SE(test_se), .CK(
        clk), .RN(n4457), .Q(RData2[29]), .QN(n82) );
  SDFFRXL \RData2_reg[28]  ( .D(next_RData2[28]), .SI(n63), .SE(test_se), .CK(
        clk), .RN(n4457), .Q(RData2[28]), .QN(n81) );
  SDFFRXL \RData1_reg[26]  ( .D(next_RData1[26]), .SI(n49), .SE(test_se), .CK(
        clk), .RN(n4454), .Q(RData1[26]), .QN(n80) );
  SDFFRXL \RData1_reg[23]  ( .D(next_RData1[23]), .SI(n48), .SE(test_se), .CK(
        clk), .RN(n4455), .Q(RData1[23]), .QN(n79) );
  SDFFRXL \RData1_reg[21]  ( .D(next_RData1[21]), .SI(n47), .SE(test_se), .CK(
        clk), .RN(n4455), .Q(RData1[21]), .QN(n78) );
  SDFFRXL \RData1_reg[19]  ( .D(next_RData1[19]), .SI(n75), .SE(test_se), .CK(
        clk), .RN(n4455), .Q(RData1[19]), .QN(n77) );
  SDFFRXL \RData1_reg[18]  ( .D(next_RData1[18]), .SI(n74), .SE(test_se), .CK(
        clk), .RN(n4455), .Q(RData1[18]), .QN(n75) );
  SDFFRXL \RData1_reg[17]  ( .D(next_RData1[17]), .SI(n72), .SE(test_se), .CK(
        clk), .RN(n4455), .Q(RData1[17]), .QN(n74) );
  SDFFRXL \RData1_reg[16]  ( .D(next_RData1[16]), .SI(n71), .SE(test_se), .CK(
        clk), .RN(n4455), .Q(RData1[16]), .QN(n72) );
  SDFFRXL \RData1_reg[15]  ( .D(next_RData1[15]), .SI(n1625), .SE(test_se), 
        .CK(clk), .RN(n4455), .Q(RData1[15]), .QN(n71) );
  SDFFRXL \RData1_reg[13]  ( .D(next_RData1[13]), .SI(n1627), .SE(test_se), 
        .CK(clk), .RN(n4456), .Q(RData1[13]), .QN(n70) );
  SDFFRXL \RData1_reg[5]  ( .D(next_RData1[5]), .SI(n1631), .SE(test_se), .CK(
        clk), .RN(n4456), .Q(RData1[5]), .QN(n69) );
  SDFFRXL \RData1_reg[2]  ( .D(next_RData1[2]), .SI(n40), .SE(test_se), .CK(
        clk), .RN(n4456), .Q(RData1[2]), .QN(n68) );
  SDFFRXL \RData2_reg[31]  ( .D(next_RData2[31]), .SI(n64), .SE(test_se), .CK(
        clk), .RN(n4457), .Q(RData2[31]), .QN(n67) );
  SDFFRXL \RData2_reg[30]  ( .D(next_RData2[30]), .SI(n82), .SE(test_se), .CK(
        clk), .RN(n4457), .Q(RData2[30]), .QN(n64) );
  SDFFRXL \RData2_reg[27]  ( .D(next_RData2[27]), .SI(n60), .SE(test_se), .CK(
        clk), .RN(n4457), .Q(RData2[27]), .QN(n63) );
  SDFFRXL \RData2_reg[26]  ( .D(next_RData2[26]), .SI(n1623), .SE(test_se), 
        .CK(clk), .RN(n4457), .Q(RData2[26]), .QN(n60) );
  SDFFRXL \RData2_reg[23]  ( .D(next_RData2[23]), .SI(n58), .SE(test_se), .CK(
        clk), .RN(n4457), .Q(RData2[23]), .QN(n59) );
  SDFFRXL \RData2_reg[22]  ( .D(next_RData2[22]), .SI(n56), .SE(test_se), .CK(
        clk), .RN(n4457), .Q(RData2[22]), .QN(n58) );
  SDFFRXL \RData2_reg[21]  ( .D(next_RData2[21]), .SI(n55), .SE(test_se), .CK(
        clk), .RN(n4458), .Q(RData2[21]), .QN(n56) );
  SDFFRXL \RData2_reg[20]  ( .D(next_RData2[20]), .SI(n52), .SE(test_se), .CK(
        clk), .RN(n4458), .Q(RData2[20]), .QN(n55) );
  SDFFRXL \RData2_reg[19]  ( .D(next_RData2[19]), .SI(n51), .SE(test_se), .CK(
        clk), .RN(n4458), .Q(RData2[19]), .QN(n52) );
  SDFFRXL \RData2_reg[18]  ( .D(next_RData2[18]), .SI(n50), .SE(test_se), .CK(
        clk), .RN(n4458), .Q(RData2[18]), .QN(n51) );
  SDFFRXL \RData2_reg[17]  ( .D(next_RData2[17]), .SI(n1667), .SE(test_se), 
        .CK(clk), .RN(n4458), .Q(RData2[17]), .QN(n50) );
  SDFFRXL \RData1_reg[25]  ( .D(next_RData1[25]), .SI(n42), .SE(test_se), .CK(
        clk), .RN(n4455), .Q(RData1[25]), .QN(n49) );
  SDFFRXL \RData1_reg[22]  ( .D(next_RData1[22]), .SI(n78), .SE(test_se), .CK(
        clk), .RN(n4455), .Q(RData1[22]), .QN(n48) );
  SDFFRXL \RData1_reg[20]  ( .D(next_RData1[20]), .SI(n77), .SE(test_se), .CK(
        clk), .RN(n4455), .Q(RData1[20]), .QN(n47) );
  SDFFRXL \RData1_reg[11]  ( .D(next_RData1[11]), .SI(n1629), .SE(test_se), 
        .CK(clk), .RN(n4456), .Q(RData1[11]), .QN(n46) );
  SDFFRXL \RData1_reg[9]  ( .D(next_RData1[9]), .SI(n1633), .SE(test_se), .CK(
        clk), .RN(n4456), .Q(RData1[9]), .QN(n45) );
  SDFFRXL \RData1_reg[7]  ( .D(next_RData1[7]), .SI(n43), .SE(test_se), .CK(
        clk), .RN(n4456), .Q(RData1[7]), .QN(n44) );
  SDFFRXL \RData1_reg[6]  ( .D(next_RData1[6]), .SI(n69), .SE(test_se), .CK(
        clk), .RN(n4456), .Q(RData1[6]), .QN(n43) );
  SDFFRXL \RData1_reg[24]  ( .D(next_RData1[24]), .SI(n79), .SE(test_se), .CK(
        clk), .RN(n4455), .Q(RData1[24]), .QN(n42) );
  SDFFRXL \RData1_reg[3]  ( .D(next_RData1[3]), .SI(n68), .SE(test_se), .CK(
        clk), .RN(n4456), .Q(RData1[3]), .QN(n41) );
  SDFFRXL \RData1_reg[1]  ( .D(next_RData1[1]), .SI(n1635), .SE(test_se), .CK(
        clk), .RN(n4457), .Q(RData1[1]), .QN(n40) );
  SDFFNSRXL \regfile_reg[3][2]  ( .D(n1746), .SI(n1547), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4514), .Q(\regfile[3][2] ), .QN(n1546) );
  SDFFRXL \Immediate_SE_reg[5]  ( .D(n146), .SI(n625), .SE(test_se), .CK(clk), 
        .RN(n4462), .Q(n1947), .QN(n626) );
  SDFFRXL \Immediate_SE_reg[2]  ( .D(n143), .SI(n612), .SE(test_se), .CK(clk), 
        .RN(n4462), .Q(n1949), .QN(n39) );
  SDFFNSRXL \regfile_reg[3][6]  ( .D(n1754), .SI(n1543), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4514), .Q(\regfile[3][6] ), .QN(n1542) );
  SDFFNSRXL \regfile_reg[3][17]  ( .D(n1776), .SI(n1532), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4513), .Q(\regfile[3][17] ), .QN(n1531) );
  SDFFNSRXL \regfile_reg[3][16]  ( .D(n1774), .SI(n1533), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4513), .Q(\regfile[3][16] ), .QN(n1532) );
  SDFFRXL \RegisterRs_reg[1]  ( .D(n3622), .SI(n648), .SE(test_se), .CK(clk), 
        .RN(n4450), .Q(RegisterRs[1]), .QN(n649) );
  SDFFNSRXL \regfile_reg[3][10]  ( .D(n1762), .SI(n1539), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4513), .Q(n88), .QN(n1538) );
  SDFFNSRXL \regfile_reg[2][29]  ( .D(n1736), .SI(n4570), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4514), .Q(n4571), .QN(n1551) );
  SDFFNSRXL \regfile_reg[2][28]  ( .D(n1734), .SI(n4569), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4514), .Q(n4570), .QN(n1552) );
  SDFFNSRXL \regfile_reg[2][26]  ( .D(n1730), .SI(n4567), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4514), .Q(n4568), .QN(n1554) );
  SDFFNSRXL \regfile_reg[2][31]  ( .D(n1740), .SI(n4572), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4514), .Q(n4573), .QN(n1549) );
  SDFFNSRXL \regfile_reg[2][30]  ( .D(n1738), .SI(n4571), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4514), .Q(n4572), .QN(n1550) );
  SDFFNSRXL \regfile_reg[2][27]  ( .D(n1732), .SI(n4568), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4514), .Q(n4569), .QN(n1553) );
  SDFFNSRXL \regfile_reg[2][9]  ( .D(n1696), .SI(n4550), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4515), .Q(n4551), .QN(n1571) );
  SDFFNSRXL \regfile_reg[2][25]  ( .D(n1728), .SI(n4566), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4514), .Q(n4567), .QN(n1555) );
  SDFFNSRXL \regfile_reg[2][10]  ( .D(n1698), .SI(n4551), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4515), .Q(n4552), .QN(n1570) );
  SDFFNSRXL \regfile_reg[2][7]  ( .D(n1692), .SI(n4548), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4515), .Q(n4549), .QN(n1573) );
  SDFFNSRXL \regfile_reg[2][6]  ( .D(n1690), .SI(n4547), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4515), .Q(n4548), .QN(n1574) );
  SDFFNSRXL \regfile_reg[2][5]  ( .D(n1688), .SI(n4546), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4515), .Q(n4547), .QN(n1575) );
  SDFFNSRXL \regfile_reg[2][2]  ( .D(n1682), .SI(n4543), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4516), .Q(n4544), .QN(n1578) );
  SDFFNSRXL \regfile_reg[2][15]  ( .D(n1708), .SI(n4556), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4515), .Q(n4557), .QN(n1565) );
  SDFFNSRXL \regfile_reg[2][12]  ( .D(n1702), .SI(n4553), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4515), .Q(n4554), .QN(n1568) );
  SDFFNSRXL \regfile_reg[2][8]  ( .D(n1694), .SI(n4549), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4515), .Q(n4550), .QN(n1572) );
  SDFFNSRXL \regfile_reg[2][24]  ( .D(n1726), .SI(n4565), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4514), .Q(n4566), .QN(n1556) );
  SDFFNSRXL \regfile_reg[2][14]  ( .D(n1706), .SI(n4555), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4515), .Q(n4556), .QN(n1566) );
  SDFFNSRXL \regfile_reg[2][4]  ( .D(n1686), .SI(n4545), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4515), .Q(n4546), .QN(n1576) );
  SDFFNSRXL \regfile_reg[2][1]  ( .D(n1680), .SI(n4542), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4516), .Q(n4543), .QN(n1579) );
  SDFFNSRXL \regfile_reg[2][3]  ( .D(n1684), .SI(n4544), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4516), .Q(n4545), .QN(n1577) );
  SDFFNSRXL \regfile_reg[2][23]  ( .D(n1724), .SI(n4564), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4514), .Q(n4565), .QN(n1557) );
  SDFFNSRXL \regfile_reg[2][22]  ( .D(n1722), .SI(n4563), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4514), .Q(n4564), .QN(n1558) );
  SDFFNSRXL \regfile_reg[2][21]  ( .D(n1720), .SI(n4562), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4515), .Q(n4563), .QN(n1559) );
  SDFFNSRXL \regfile_reg[2][20]  ( .D(n1718), .SI(n4561), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4515), .Q(n4562), .QN(n1560) );
  SDFFNSRXL \regfile_reg[2][19]  ( .D(n1716), .SI(n4560), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4515), .Q(n4561), .QN(n1561) );
  SDFFNSRXL \regfile_reg[2][18]  ( .D(n1714), .SI(n4559), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4515), .Q(n4560), .QN(n1562) );
  SDFFNSRXL \regfile_reg[2][17]  ( .D(n1712), .SI(n4558), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4515), .Q(n4559), .QN(n1563) );
  SDFFNSRXL \regfile_reg[2][16]  ( .D(n1710), .SI(n4557), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4515), .Q(n4558), .QN(n1564) );
  SDFFNSRXL \regfile_reg[2][13]  ( .D(n1704), .SI(n4554), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4515), .Q(n4555), .QN(n1567) );
  SDFFNSRXL \regfile_reg[2][11]  ( .D(n1700), .SI(n4552), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4515), .Q(n4553), .QN(n1569) );
  SDFFNSRXL \regfile_reg[2][0]  ( .D(n1678), .SI(n1581), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4516), .Q(n4542), .QN(n1580) );
  SDFFRXL \PCBuffer_reg[31]  ( .D(n3587), .SI(n17), .SE(test_se), .CK(clk), 
        .RN(rst), .Q(n4639), .QN(n3626) );
  SDFFRXL \EX_reg[0]  ( .D(n3605), .SI(test_si2), .SE(test_se), .CK(clk), .RN(
        n4451), .Q(EX[0]), .QN(n38) );
  SDFFRXL \EX_reg[4]  ( .D(n3609), .SI(n640), .SE(test_se), .CK(clk), .RN(
        n4451), .Q(n1941), .QN(n37) );
  SDFFRXL \RegisterRs_reg[0]  ( .D(n3621), .SI(n635), .SE(test_se), .CK(clk), 
        .RN(n4450), .Q(RegisterRs[0]), .QN(n648) );
  SDFFRXL \RegisterRs_reg[3]  ( .D(n3624), .SI(n650), .SE(test_se), .CK(clk), 
        .RN(n4450), .Q(RegisterRs[3]), .QN(n651) );
  SDFFRXL \RegisterRs_reg[2]  ( .D(n3623), .SI(n649), .SE(test_se), .CK(clk), 
        .RN(n4450), .Q(RegisterRs[2]), .QN(n650) );
  SDFFRXL \RegisterRt_reg[1]  ( .D(n3617), .SI(n643), .SE(test_se), .CK(clk), 
        .RN(n4450), .Q(n1959), .QN(n644) );
  SDFFRXL \RegisterRt_reg[4]  ( .D(n3620), .SI(n646), .SE(test_se), .CK(clk), 
        .RN(n4450), .Q(n1953), .QN(n647) );
  SDFFRXL \RegisterRt_reg[2]  ( .D(n3618), .SI(n644), .SE(test_se), .CK(clk), 
        .RN(n4450), .Q(n1957), .QN(n645) );
  SDFFRXL \RegisterRt_reg[3]  ( .D(n3619), .SI(n645), .SE(test_se), .CK(clk), 
        .RN(n4450), .Q(n1955), .QN(n646) );
  SDFFRXL \RegisterRt_reg[0]  ( .D(n3616), .SI(n652), .SE(test_se), .CK(clk), 
        .RN(n4450), .Q(n1961), .QN(n643) );
  SDFFRXL \Immediate_SE_reg[20]  ( .D(next_Immediate_SE[20]), .SI(n611), .SE(
        test_se), .CK(clk), .RN(n4460), .Q(Immediate_SE[20]), .QN(n613) );
  SDFFRXL \Immediate_SE_reg[25]  ( .D(next_Immediate_SE[25]), .SI(n617), .SE(
        test_se), .CK(clk), .RN(n4460), .Q(Immediate_SE[25]), .QN(n618) );
  SDFFRXL \Immediate_SE_reg[24]  ( .D(next_Immediate_SE[24]), .SI(n616), .SE(
        test_se), .CK(clk), .RN(n4460), .Q(Immediate_SE[24]), .QN(n617) );
  SDFFNSRXL \regfile_reg[3][7]  ( .D(n1756), .SI(n1542), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4514), .Q(n89), .QN(n1541) );
  SDFFNSRXL \regfile_reg[3][4]  ( .D(n1750), .SI(\regfile[3][3] ), .SE(test_se), .CKN(clk), .SN(1'b1), .RN(n4514), .Q(n90), .QN(n1544) );
  SDFFNSRXL \regfile_reg[3][3]  ( .D(n1748), .SI(n1546), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4514), .Q(\regfile[3][3] ), .QN(n1545) );
  SDFFNSRXL \regfile_reg[3][23]  ( .D(n1788), .SI(n1526), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4513), .Q(n87), .QN(n1525) );
  SDFFNSRXL \regfile_reg[3][20]  ( .D(n1782), .SI(n1529), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4513), .Q(n85), .QN(n1528) );
  SDFFNSRXL \regfile_reg[3][19]  ( .D(n1780), .SI(n1530), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4513), .Q(n94), .QN(n1529) );
  SDFFNSRXL \regfile_reg[3][18]  ( .D(n1778), .SI(n1531), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4513), .Q(n91), .QN(n1530) );
  SDFFNSRXL \regfile_reg[3][0]  ( .D(n1742), .SI(n4573), .SE(test_se), .CKN(
        clk), .SN(1'b1), .RN(n4514), .Q(n92), .QN(n1548) );
  INVXL U1 ( .A(\regfile[1][0] ), .Y(n1757) );
  INVXL U2 ( .A(\regfile[1][2] ), .Y(n1759) );
  INVXL U3 ( .A(\regfile[1][5] ), .Y(n1763) );
  INVXL U4 ( .A(\regfile[1][8] ), .Y(n1765) );
  INVXL U10 ( .A(\regfile[1][24] ), .Y(n1767) );
  INVXL U13 ( .A(\regfile[1][3] ), .Y(n1769) );
  INVXL U31 ( .A(\regfile[1][4] ), .Y(n1771) );
  INVXL U32 ( .A(\regfile[1][9] ), .Y(n1773) );
  INVXL U34 ( .A(\regfile[1][19] ), .Y(n1775) );
  INVXL U36 ( .A(\regfile[1][30] ), .Y(n1783) );
  MXI2X4 U37 ( .A(n516), .B(n1553), .S0(n1857), .Y(n519) );
  NOR2BX4 U39 ( .AN(n1601), .B(n4270), .Y(n4199) );
  CLKAND2X12 U40 ( .A(n4424), .B(n1588), .Y(n4134) );
  AOI221X4 U41 ( .A0(n1891), .A1(EX_RegWriteData[3]), .B0(next_RData1[3]), 
        .B1(n1889), .C0(n1789), .Y(n1785) );
  CLKINVX20 U42 ( .A(n1785), .Y(n4948) );
  CLKINVX20 U47 ( .A(n4940), .Y(n1789) );
  MXI2X4 U88 ( .A(n4162), .B(n1562), .S0(n1863), .Y(n4165) );
  NOR2BX4 U89 ( .AN(n1596), .B(n3742), .Y(n630) );
  NAND4X8 U90 ( .A(n1791), .B(n4930), .C(n4929), .D(n4928), .Y(n4979) );
  CLKXOR2X8 U91 ( .A(n1801), .B(n4899), .Y(n1791) );
  CLKBUFX20 U92 ( .A(n4643), .Y(n1793) );
  CLKAND2X12 U93 ( .A(Branch), .B(equal), .Y(n1795) );
  AOI221X4 U94 ( .A0(n1891), .A1(EX_RegWriteData[14]), .B0(next_RData1[14]), 
        .B1(n1889), .C0(n1799), .Y(n1797) );
  CLKINVX20 U95 ( .A(n1797), .Y(n4821) );
  CLKINVX20 U96 ( .A(n4813), .Y(n1799) );
  CLKAND2X12 U97 ( .A(n4424), .B(n1612), .Y(n4254) );
  AND3X8 U98 ( .A(n95), .B(n96), .C(n4892), .Y(n1801) );
  CLKAND2X12 U99 ( .A(n1803), .B(n1610), .Y(n3719) );
  CLKINVX20 U100 ( .A(n3746), .Y(n1803) );
  CLKMX2X6 U101 ( .A(n1807), .B(n1805), .S0(n4257), .Y(N148) );
  MXI4X4 U102 ( .A(n4092), .B(n4090), .C(n4091), .D(n4089), .S0(N25), .S1(
        n4265), .Y(n1805) );
  MXI4X4 U103 ( .A(n4096), .B(n4094), .C(n4095), .D(n4093), .S0(N25), .S1(
        n4265), .Y(n1807) );
  CLKAND2X12 U104 ( .A(n1603), .B(n1809), .Y(n4209) );
  CLKINVX20 U105 ( .A(n4280), .Y(n1809) );
  OR2X8 U106 ( .A(n4244), .B(n4243), .Y(n1811) );
  CLKINVX20 U107 ( .A(n1811), .Y(n4246) );
  AOI221X4 U108 ( .A0(n1891), .A1(EX_RegWriteData[4]), .B0(next_RData1[4]), 
        .B1(n1889), .C0(n1815), .Y(n1813) );
  CLKINVX20 U109 ( .A(n1813), .Y(n4918) );
  CLKINVX20 U110 ( .A(n4910), .Y(n1815) );
  MXI2X4 U111 ( .A(n4172), .B(n1564), .S0(n1863), .Y(n4175) );
  MXI2X4 U112 ( .A(n1741), .B(n1571), .S0(n1857), .Y(n1755) );
  AOI221X4 U113 ( .A0(n1891), .A1(EX_RegWriteData[21]), .B0(next_RData1[21]), 
        .B1(n1889), .C0(n1819), .Y(n1817) );
  CLKINVX20 U114 ( .A(n1817), .Y(n4764) );
  CLKINVX20 U115 ( .A(n4756), .Y(n1819) );
  MXI2X4 U116 ( .A(n3808), .B(n3807), .S0(n4428), .Y(N164) );
  CLKMX2X6 U117 ( .A(n1823), .B(n1821), .S0(n4257), .Y(N158) );
  MXI4X4 U118 ( .A(n4012), .B(n4010), .C(n4011), .D(n4009), .S0(n4261), .S1(
        n4264), .Y(n1821) );
  MXI4X4 U119 ( .A(n4016), .B(n4014), .C(n4015), .D(n4013), .S0(n4261), .S1(
        n4264), .Y(n1823) );
  CLKAND2X12 U120 ( .A(n4431), .B(n1604), .Y(n1781) );
  CLKAND2X12 U121 ( .A(n1582), .B(n1825), .Y(n503) );
  CLKINVX20 U122 ( .A(n3748), .Y(n1825) );
  MXI2X4 U123 ( .A(n4217), .B(n1573), .S0(n1863), .Y(n4220) );
  MXI2X4 U124 ( .A(n4187), .B(n1567), .S0(n1863), .Y(n4190) );
  MXI2X4 U125 ( .A(n4132), .B(n1556), .S0(n1863), .Y(n4135) );
  AOI221X4 U126 ( .A0(n1891), .A1(EX_RegWriteData[1]), .B0(next_RData1[1]), 
        .B1(n1889), .C0(n1829), .Y(n1827) );
  CLKINVX20 U127 ( .A(n1827), .Y(n4974) );
  CLKINVX20 U128 ( .A(n4960), .Y(n1829) );
  MXI2X4 U174 ( .A(n3727), .B(n1580), .S0(n1857), .Y(n3730) );
  MXI2X4 U236 ( .A(n3822), .B(n3821), .S0(n1893), .Y(N157) );
  CLKAND2X12 U241 ( .A(n1593), .B(n1831), .Y(n4159) );
  CLKINVX20 U242 ( .A(n4268), .Y(n1831) );
  MXI2X4 U249 ( .A(n4252), .B(n1580), .S0(n1863), .Y(n4255) );
  CLKAND2X12 U268 ( .A(n1609), .B(n1833), .Y(n4239) );
  CLKINVX20 U271 ( .A(n4270), .Y(n1833) );
  MXI2X4 U279 ( .A(n3717), .B(n1578), .S0(n1857), .Y(n3720) );
  MXI2X4 U280 ( .A(n3830), .B(n3829), .S0(n1893), .Y(N153) );
  MXI2X4 U282 ( .A(n4197), .B(n1569), .S0(n1863), .Y(n4200) );
  MXI2X4 U283 ( .A(n628), .B(n1564), .S0(n1857), .Y(n1677) );
  CLKAND2X12 U284 ( .A(n1608), .B(n1835), .Y(n4234) );
  CLKINVX20 U288 ( .A(n4269), .Y(n1835) );
  MXI2X4 U293 ( .A(n3790), .B(n3789), .S0(n1893), .Y(N173) );
  MXI2X4 U303 ( .A(n3780), .B(n3779), .S0(n1893), .Y(N178) );
  CLKAND2X12 U343 ( .A(n4424), .B(n1607), .Y(n4229) );
  MXI2X4 U534 ( .A(n4242), .B(n1578), .S0(n1863), .Y(n4245) );
  CLKMX2X6 U659 ( .A(n1839), .B(n1837), .S0(n3732), .Y(N142) );
  MXI4X4 U724 ( .A(n283), .B(n281), .C(n282), .D(n280), .S0(n3734), .S1(n3738), 
        .Y(n1837) );
  MXI4X4 U879 ( .A(n287), .B(n285), .C(n286), .D(n284), .S0(n3734), .S1(n3738), 
        .Y(n1839) );
  MXI2X4 U883 ( .A(n3832), .B(n3831), .S0(n1893), .Y(N152) );
  MXI2X4 U884 ( .A(n3812), .B(n3811), .S0(n1893), .Y(N162) );
  CLKMX2X6 U885 ( .A(n1843), .B(n1841), .S0(N26), .Y(N167) );
  MXI4X4 U886 ( .A(n3940), .B(n3938), .C(n3939), .D(n3937), .S0(n4258), .S1(
        n4262), .Y(n1841) );
  MXI4X4 U887 ( .A(n3944), .B(n3942), .C(n3943), .D(n3941), .S0(n4258), .S1(
        N24), .Y(n1843) );
  MXI2X4 U894 ( .A(n3697), .B(n1574), .S0(n1857), .Y(n3700) );
  CLKMX2X6 U895 ( .A(n1847), .B(n1845), .S0(n4257), .Y(N159) );
  MXI4X4 U906 ( .A(n4004), .B(n4002), .C(n4003), .D(n4001), .S0(n4261), .S1(
        n4264), .Y(n1845) );
  MXI4X4 U916 ( .A(n4008), .B(n4006), .C(n4007), .D(n4005), .S0(n4261), .S1(
        n4264), .Y(n1847) );
  MXI2X4 U919 ( .A(n4127), .B(n1555), .S0(n1863), .Y(n4130) );
  MXI2X4 U920 ( .A(n4212), .B(n1572), .S0(n1863), .Y(n4215) );
  AOI221X4 U929 ( .A0(n1891), .A1(EX_RegWriteData[20]), .B0(next_RData1[20]), 
        .B1(n1889), .C0(n1851), .Y(n1849) );
  CLKINVX20 U930 ( .A(n1849), .Y(n4755) );
  CLKINVX20 U931 ( .A(n4747), .Y(n1851) );
  MXI2X4 U946 ( .A(n1701), .B(n1567), .S0(n1857), .Y(n1707) );
  MXI2X4 U997 ( .A(n1777), .B(n1572), .S0(n1857), .Y(n1787) );
  MXI2X4 U998 ( .A(n506), .B(n1551), .S0(n1857), .Y(n509) );
  MXI2X4 U1043 ( .A(n4157), .B(n1561), .S0(n1863), .Y(n4160) );
  AOI221X4 U1051 ( .A0(EX_RegWriteData[19]), .A1(n1891), .B0(next_RData1[19]), 
        .B1(n1889), .C0(n1855), .Y(n1853) );
  CLKINVX20 U1083 ( .A(n1853), .Y(n4786) );
  OAI22X4 U1087 ( .A0(n4781), .A1(n4403), .B0(n4780), .B1(n4400), .Y(n1855) );
  MXI2X4 U1127 ( .A(n4207), .B(n1571), .S0(n1863), .Y(n4210) );
  MXI2X4 U1143 ( .A(n3834), .B(n3833), .S0(n1893), .Y(N151) );
  MXI2X4 U1263 ( .A(n4107), .B(n1551), .S0(n1863), .Y(n4110) );
  MXI2X4 U1266 ( .A(n521), .B(n1554), .S0(n1857), .Y(n524) );
  CLKINVX20 U1273 ( .A(n3774), .Y(n1857) );
  AOI221X4 U1274 ( .A0(n1891), .A1(EX_RegWriteData[23]), .B0(next_RData1[23]), 
        .B1(n1889), .C0(n1861), .Y(n1859) );
  CLKINVX20 U1276 ( .A(n1859), .Y(n4746) );
  OAI22X4 U1277 ( .A0(n4402), .A1(n4741), .B0(n4401), .B1(n4740), .Y(n1861) );
  MXI2X4 U1279 ( .A(n4232), .B(n1576), .S0(n1863), .Y(n4235) );
  CLKINVX20 U1281 ( .A(n4298), .Y(n1863) );
  AOI221X4 U1283 ( .A0(n1891), .A1(EX_RegWriteData[22]), .B0(next_RData1[22]), 
        .B1(n1889), .C0(n1867), .Y(n1865) );
  CLKINVX20 U1284 ( .A(n1865), .Y(n4737) );
  OAI22X4 U1285 ( .A0(n4403), .A1(n4732), .B0(n4401), .B1(n4731), .Y(n1867) );
  AOI221X4 U1286 ( .A0(n1891), .A1(EX_RegWriteData[17]), .B0(next_RData1[17]), 
        .B1(n1889), .C0(n1871), .Y(n1869) );
  CLKINVX20 U1287 ( .A(n1869), .Y(n4804) );
  OAI22X4 U1290 ( .A0(n4402), .A1(n4799), .B0(n4401), .B1(n4798), .Y(n1871) );
  MXI2X4 U1292 ( .A(n4222), .B(n1574), .S0(n4423), .Y(n4225) );
  MXI2X4 U1294 ( .A(n4227), .B(n1575), .S0(n4423), .Y(n4230) );
  AOI221X4 U1297 ( .A0(n1891), .A1(EX_RegWriteData[12]), .B0(next_RData1[12]), 
        .B1(n1889), .C0(n1875), .Y(n1873) );
  CLKINVX20 U1299 ( .A(n1873), .Y(n4839) );
  CLKINVX20 U1300 ( .A(n4831), .Y(n1875) );
  MXI2X4 U1337 ( .A(n3838), .B(n3837), .S0(n1893), .Y(N149) );
  AOI221X4 U1341 ( .A0(n1891), .A1(EX_RegWriteData[28]), .B0(next_RData1[28]), 
        .B1(n1889), .C0(n1879), .Y(n1877) );
  CLKINVX20 U1349 ( .A(n1877), .Y(n4675) );
  OAI22X4 U1363 ( .A0(n4403), .A1(n4670), .B0(n4400), .B1(n4669), .Y(n1879) );
  CLKMX2X6 U1369 ( .A(n1883), .B(n1881), .S0(N26), .Y(N169) );
  MXI4X4 U1370 ( .A(n3924), .B(n3922), .C(n3923), .D(n3921), .S0(n4258), .S1(
        n4263), .Y(n1881) );
  MXI4X4 U1378 ( .A(n3928), .B(n3926), .C(n3927), .D(n3925), .S0(n4426), .S1(
        n4265), .Y(n1883) );
  AOI221X4 U1382 ( .A0(n1891), .A1(EX_RegWriteData[7]), .B0(next_RData1[7]), 
        .B1(n1889), .C0(n1887), .Y(n1885) );
  CLKINVX20 U1386 ( .A(n1885), .Y(n4909) );
  CLKINVX20 U1390 ( .A(n4901), .Y(n1887) );
  CLKINVX20 U1394 ( .A(n4404), .Y(n1889) );
  CLKINVX20 U1398 ( .A(n4406), .Y(n1891) );
  MXI2X4 U1405 ( .A(n3806), .B(n3805), .S0(n1893), .Y(N165) );
  CLKINVX20 U1413 ( .A(N26), .Y(n1893) );
  MXI2X4 U1425 ( .A(n531), .B(n1556), .S0(n4430), .Y(n534) );
  MXI2X4 U1433 ( .A(n501), .B(n1550), .S0(n4430), .Y(n504) );
  CLKBUFX20 U1437 ( .A(n1538), .Y(n1895) );
  CLKAND2X12 U1457 ( .A(n4268), .B(n1895), .Y(n4202) );
  INVXL U1465 ( .A(n3658), .Y(n1897) );
  INVXL U1473 ( .A(n1897), .Y(n1899) );
  INVXL U1488 ( .A(n1897), .Y(n1901) );
  CLKBUFX2 U1496 ( .A(n1915), .Y(Immediate_SE[2]) );
  CLKBUFX2 U1500 ( .A(n1951), .Y(Immediate_SE[1]) );
  CLKBUFX2 U1516 ( .A(n1945), .Y(EX[1]) );
  CLKBUFX2 U1528 ( .A(n1943), .Y(EX[2]) );
  INVXL U1560 ( .A(n1949), .Y(n1911) );
  INVXL U1564 ( .A(n1911), .Y(n1913) );
  INVXL U1568 ( .A(n1911), .Y(n1915) );
  CLKBUFX2 U1576 ( .A(n1957), .Y(RegisterRt[2]) );
  CLKBUFX2 U1580 ( .A(n1959), .Y(RegisterRt[1]) );
  CLKBUFX2 U1596 ( .A(n1955), .Y(RegisterRt[3]) );
  CLKBUFX2 U1604 ( .A(n1961), .Y(RegisterRt[0]) );
  CLKBUFX2 U1612 ( .A(n1953), .Y(RegisterRt[4]) );
  CLKBUFX2 U1685 ( .A(n1931), .Y(Immediate_SE[5]) );
  INVXL U1686 ( .A(n1947), .Y(n1929) );
  INVXL U1687 ( .A(n1929), .Y(n1931) );
  CLKBUFX2 U1688 ( .A(n1937), .Y(EX[4]) );
  INVXL U1689 ( .A(n1941), .Y(n1935) );
  INVXL U1690 ( .A(n1935), .Y(n1937) );
  INVXL U1691 ( .A(n1935), .Y(n1939) );
endmodule


module InstructionFetch_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32;

  AND2X2 U1 ( .A(A[30]), .B(n28), .Y(n1) );
  AND2X2 U2 ( .A(A[29]), .B(n27), .Y(n28) );
  XOR2X1 U3 ( .A(A[29]), .B(n27), .Y(SUM[29]) );
  XOR2X1 U4 ( .A(A[30]), .B(n28), .Y(SUM[30]) );
  XOR2X1 U5 ( .A(A[31]), .B(n1), .Y(SUM[31]) );
  AND2XL U6 ( .A(A[13]), .B(n12), .Y(n13) );
  AND2XL U7 ( .A(A[15]), .B(n14), .Y(n15) );
  AND2XL U8 ( .A(A[14]), .B(n13), .Y(n14) );
  AND2XL U9 ( .A(A[16]), .B(n15), .Y(n16) );
  AND2XL U10 ( .A(A[17]), .B(n16), .Y(n17) );
  AND2XL U11 ( .A(A[18]), .B(n17), .Y(n18) );
  AND2XL U12 ( .A(A[19]), .B(n18), .Y(n19) );
  AND2XL U13 ( .A(A[20]), .B(n19), .Y(n20) );
  AND2XL U14 ( .A(A[21]), .B(n20), .Y(n21) );
  AND2XL U15 ( .A(A[22]), .B(n21), .Y(n22) );
  AND2XL U16 ( .A(n30), .B(n29), .Y(n23) );
  AND2XL U18 ( .A(A[25]), .B(n24), .Y(n2) );
  AND2XL U19 ( .A(A[27]), .B(n25), .Y(n26) );
  AND2XL U20 ( .A(A[26]), .B(n2), .Y(n25) );
  AND2XL U21 ( .A(A[28]), .B(n26), .Y(n27) );
  AND2XL U22 ( .A(A[3]), .B(A[2]), .Y(n3) );
  AND2XL U23 ( .A(A[4]), .B(n3), .Y(n4) );
  AND2XL U24 ( .A(A[5]), .B(n4), .Y(n5) );
  AND2XL U25 ( .A(A[6]), .B(n5), .Y(n6) );
  AND2XL U26 ( .A(A[7]), .B(n6), .Y(n7) );
  AND2XL U27 ( .A(A[8]), .B(n7), .Y(n8) );
  AND2XL U28 ( .A(A[9]), .B(n8), .Y(n9) );
  AND2XL U29 ( .A(A[10]), .B(n9), .Y(n10) );
  AND2XL U30 ( .A(A[11]), .B(n10), .Y(n11) );
  AND2XL U31 ( .A(A[12]), .B(n11), .Y(n12) );
  XOR2XL U32 ( .A(A[28]), .B(n26), .Y(SUM[28]) );
  INVXL U33 ( .A(A[2]), .Y(SUM[2]) );
  XOR2XL U34 ( .A(A[14]), .B(n13), .Y(SUM[14]) );
  XOR2XL U35 ( .A(A[3]), .B(A[2]), .Y(SUM[3]) );
  XOR2XL U36 ( .A(A[4]), .B(n3), .Y(SUM[4]) );
  XOR2XL U37 ( .A(A[6]), .B(n5), .Y(SUM[6]) );
  XOR2XL U38 ( .A(A[7]), .B(n6), .Y(SUM[7]) );
  XOR2XL U39 ( .A(A[8]), .B(n7), .Y(SUM[8]) );
  XOR2XL U40 ( .A(A[9]), .B(n8), .Y(SUM[9]) );
  XOR2XL U41 ( .A(A[10]), .B(n9), .Y(SUM[10]) );
  XOR2XL U42 ( .A(A[11]), .B(n10), .Y(SUM[11]) );
  XOR2XL U43 ( .A(A[12]), .B(n11), .Y(SUM[12]) );
  XOR2XL U44 ( .A(A[13]), .B(n12), .Y(SUM[13]) );
  XOR2XL U45 ( .A(A[15]), .B(n14), .Y(SUM[15]) );
  XOR2XL U46 ( .A(A[16]), .B(n15), .Y(SUM[16]) );
  XOR2XL U47 ( .A(A[17]), .B(n16), .Y(SUM[17]) );
  XOR2XL U48 ( .A(A[18]), .B(n17), .Y(SUM[18]) );
  XOR2XL U49 ( .A(A[19]), .B(n18), .Y(SUM[19]) );
  XOR2XL U50 ( .A(A[20]), .B(n19), .Y(SUM[20]) );
  XOR2XL U51 ( .A(A[21]), .B(n20), .Y(SUM[21]) );
  XOR2XL U52 ( .A(A[22]), .B(n21), .Y(SUM[22]) );
  XOR2XL U53 ( .A(n30), .B(n29), .Y(SUM[23]) );
  XOR2XL U54 ( .A(A[24]), .B(n23), .Y(SUM[24]) );
  XOR2XL U55 ( .A(A[25]), .B(n24), .Y(SUM[25]) );
  XOR2XL U56 ( .A(A[26]), .B(n2), .Y(SUM[26]) );
  XOR2XL U57 ( .A(A[27]), .B(n25), .Y(SUM[27]) );
  XOR2XL U58 ( .A(A[5]), .B(n4), .Y(SUM[5]) );
  CLKBUFX2 U59 ( .A(A[1]), .Y(SUM[1]) );
  CLKBUFX2 U60 ( .A(A[0]), .Y(SUM[0]) );
  CLKBUFX2 U17 ( .A(n22), .Y(n29) );
  CLKBUFX2 U61 ( .A(A[23]), .Y(n30) );
  CLKAND2X12 U62 ( .A(n29), .B(A[24]), .Y(n31) );
  NOR2BX4 U63 ( .AN(n30), .B(n32), .Y(n24) );
  CLKINVX20 U64 ( .A(n31), .Y(n32) );
endmodule


module InstructionFetch_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  ADDFXL U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  ADDFXL U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  ADDFXL U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  ADDFXL U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  ADDFXL U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  ADDFXL U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ADDFXL U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ADDFXL U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  ADDFXL U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  ADDFX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  ADDFX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  ADDFX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  ADDFX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  ADDFX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  ADDFX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ADDFHX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  CMPR32X2 U1_25 ( .A(A[25]), .B(B[25]), .C(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  ADDFHX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  ADDFHX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  ADDFHX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  ADDFXL U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  XOR3X2 U1_31 ( .A(A[31]), .B(B[31]), .C(carry[31]), .Y(SUM[31]) );
  ADDFX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  ADDFHX2 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  ADDFHX2 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  ADDFHX2 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFHX4 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFHX2 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  ADDFHX4 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  AND2X2 U1 ( .A(B[2]), .B(A[2]), .Y(n1) );
  XOR2XL U2 ( .A(B[2]), .B(A[2]), .Y(SUM[2]) );
  CLKBUFX3 U3 ( .A(A[1]), .Y(SUM[1]) );
  CLKBUFX3 U4 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module InstructionFetch_test_1 ( clk, rst, stall, PCWrite, PCJumpJRorBranch, 
        IF_ID_Write, IF_Flush, PCadd4, Instruction, PC, read_Instruction, 
        PredictMiss, BranchTaken, PCBuffer_valid, test_si, test_so, test_se );
  input [31:0] PCJumpJRorBranch;
  output [31:0] PCadd4;
  output [31:0] Instruction;
  output [31:0] PC;
  input [31:0] read_Instruction;
  input clk, rst, stall, PCWrite, IF_ID_Write, IF_Flush, PredictMiss,
         PCBuffer_valid, test_si, test_se;
  output BranchTaken, test_so;
  wire   n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n313, n314, n315,
         n316, n317, n318, n319, n321, n322, n323, n324, n325, n326, n328,
         n329, n330, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, next_BranchTaken, N13, \state[1] , N23, N24, N25, N26,
         N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54,
         N73, N74, N109, N110, N111, N112, N113, N114, n8, n45, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n104, n105, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165,
         N164, N163, N162, N161, n2, n3, n4, n5, n6, n7, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n35, n37, n39, n41, n43, n46, n48, n50,
         n54, n102, n106, n126, n184, n186, n188, n190, n192, n196, n198, n200,
         n202, n204, n208, n210, n212, n214, n216, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n34, n36,
         n38, n40, n42, n44, n47, n49, n51, n53, n55, n103, n107, n183, n185,
         n187, n189, n191, n193, n195, n197, n199, n201, n203, n205, n207,
         n209, n211, n213, n215, n217, n311, n312, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n410, n412, n413, n415, n416, n418,
         n419, n421, n422, n424, n425, n427, n428, n430, n435, n437, n439,
         n441, n442, n444, n451, n453, n454, n456, n457, n459, n460, n462,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n582, n583, n584;
  wire   [31:0] PCBrPredict;
  wire   [29:26] PCJumpEarly;
  wire   [1:0] next_state;

  TLATX1 \next_state_reg[1]  ( .G(n232), .D(N74), .Q(next_state[1]) );
  MXI2X1 U3 ( .A(n494), .B(N54), .S0(n232), .Y(n264) );
  NAND4BBXL U4 ( .AN(read_Instruction[28]), .BN(read_Instruction[29]), .C(n308), .D(n128), .Y(n125) );
  NOR3X1 U5 ( .A(read_Instruction[1]), .B(read_Instruction[27]), .C(
        read_Instruction[26]), .Y(n127) );
  NAND2X1 U7 ( .A(n266), .B(n265), .Y(n129) );
  NAND2X1 U8 ( .A(n275), .B(n274), .Y(n132) );
  NAND2X1 U9 ( .A(n269), .B(n268), .Y(n130) );
  NAND2X1 U10 ( .A(n272), .B(n271), .Y(n131) );
  NAND2X4 U11 ( .A(n287), .B(n279), .Y(n123) );
  OAI211X1 U12 ( .A0(n240), .A1(n306), .B0(n92), .C0(n93), .Y(n152) );
  OAI211X1 U13 ( .A0(n240), .A1(n305), .B0(n90), .C0(n91), .Y(n151) );
  OAI211X1 U14 ( .A0(n240), .A1(n304), .B0(n88), .C0(n89), .Y(n150) );
  OAI211X1 U15 ( .A0(n240), .A1(n302), .B0(n84), .C0(n85), .Y(n148) );
  OAI211X1 U16 ( .A0(n240), .A1(n301), .B0(n82), .C0(n83), .Y(n147) );
  OAI211X1 U17 ( .A0(n239), .A1(n300), .B0(n80), .C0(n81), .Y(n146) );
  OAI211X1 U18 ( .A0(n239), .A1(n298), .B0(n76), .C0(n77), .Y(n144) );
  OAI211X1 U19 ( .A0(n239), .A1(n296), .B0(n72), .C0(n73), .Y(n142) );
  OAI211X1 U20 ( .A0(n239), .A1(n295), .B0(n70), .C0(n71), .Y(n141) );
  OAI211X1 U21 ( .A0(n239), .A1(n294), .B0(n68), .C0(n69), .Y(n140) );
  OAI211X1 U22 ( .A0(n239), .A1(n293), .B0(n66), .C0(n67), .Y(n139) );
  OAI211X1 U23 ( .A0(n239), .A1(n292), .B0(n64), .C0(n65), .Y(n138) );
  OAI211X1 U24 ( .A0(n239), .A1(n291), .B0(n62), .C0(n63), .Y(n137) );
  OAI211X1 U25 ( .A0(n239), .A1(n290), .B0(n60), .C0(n61), .Y(n136) );
  OAI211X1 U26 ( .A0(n239), .A1(n289), .B0(n58), .C0(n59), .Y(n135) );
  OAI211X1 U27 ( .A0(n239), .A1(n288), .B0(n56), .C0(n57), .Y(n134) );
  MX2X1 U29 ( .A(n569), .B(N43), .S0(n232), .Y(n2) );
  MX2X1 U30 ( .A(n490), .B(N26), .S0(n232), .Y(n3) );
  MX2XL U31 ( .A(n515), .B(N44), .S0(n232), .Y(n4) );
  MX2X1 U32 ( .A(n539), .B(N46), .S0(n232), .Y(n5) );
  MX2X1 U33 ( .A(n542), .B(N47), .S0(n232), .Y(n6) );
  CLKMX2X2 U34 ( .A(n509), .B(N45), .S0(n232), .Y(n7) );
  CLKMX2X2 U35 ( .A(n560), .B(N42), .S0(n232), .Y(n9) );
  CLKMX2X2 U36 ( .A(n533), .B(N40), .S0(n232), .Y(n10) );
  CLKMX2X2 U37 ( .A(n554), .B(N41), .S0(n232), .Y(n11) );
  CLKINVX1 U38 ( .A(n45), .Y(n241) );
  CLKINVX1 U39 ( .A(n259), .Y(n278) );
  CLKBUFX3 U40 ( .A(n278), .Y(n230) );
  CLKMX2X2 U41 ( .A(n536), .B(N27), .S0(n232), .Y(n14) );
  CLKMX2X2 U42 ( .A(n545), .B(N29), .S0(n232), .Y(n15) );
  CLKMX2X2 U43 ( .A(n500), .B(N50), .S0(n232), .Y(n16) );
  CLKMX2X2 U44 ( .A(n563), .B(N48), .S0(n232), .Y(n17) );
  CLKMX2X2 U45 ( .A(n512), .B(N49), .S0(n232), .Y(n18) );
  AND4X1 U46 ( .A(n256), .B(n235), .C(n257), .D(n262), .Y(n19) );
  AND4X4 U47 ( .A(n121), .B(n112), .C(n108), .D(n122), .Y(N13) );
  AND4X1 U48 ( .A(PCBuffer_valid), .B(n310), .C(read_Instruction[3]), .D(n127), 
        .Y(n20) );
  BUFX4 U49 ( .A(n115), .Y(n237) );
  CLKMX2X2 U50 ( .A(n571), .B(N30), .S0(n232), .Y(n21) );
  CLKMX2X2 U51 ( .A(n524), .B(N32), .S0(n232), .Y(n22) );
  CLKMX2X2 U52 ( .A(n527), .B(N34), .S0(n232), .Y(n23) );
  CLKMX2X2 U53 ( .A(n566), .B(N33), .S0(n232), .Y(n24) );
  CLKMX2X2 U54 ( .A(n506), .B(N31), .S0(n232), .Y(n25) );
  CLKMX2X2 U55 ( .A(n548), .B(N35), .S0(n232), .Y(n26) );
  CLKMX2X2 U56 ( .A(n575), .B(N38), .S0(n232), .Y(n27) );
  CLKMX2X2 U57 ( .A(n551), .B(N37), .S0(n232), .Y(n28) );
  CLKMX2X2 U58 ( .A(n530), .B(N36), .S0(n232), .Y(n29) );
  CLKMX2X2 U59 ( .A(n557), .B(N39), .S0(n232), .Y(n30) );
  AND2X2 U61 ( .A(n380), .B(read_Instruction[15]), .Y(n224) );
  NAND4BBXL U62 ( .AN(Instruction[26]), .BN(n584), .C(n124), .D(
        Instruction[28]), .Y(n120) );
  INVX12 U63 ( .A(n32), .Y(PC[1]) );
  INVX12 U64 ( .A(n31), .Y(PC[0]) );
  MXI2X1 U65 ( .A(n485), .B(N52), .S0(n232), .Y(n270) );
  INVX3 U67 ( .A(n117), .Y(n284) );
  MXI2X1 U68 ( .A(n503), .B(N53), .S0(n279), .Y(n267) );
  INVX12 U69 ( .A(n35), .Y(PC[31]) );
  AO21X4 U70 ( .A0(PCBrPredict[31]), .A1(n229), .B0(n260), .Y(n282) );
  INVX12 U71 ( .A(n37), .Y(PC[25]) );
  INVX12 U72 ( .A(n405), .Y(PC[27]) );
  INVX12 U73 ( .A(n399), .Y(PC[26]) );
  INVX12 U74 ( .A(n402), .Y(PC[28]) );
  INVX12 U75 ( .A(n396), .Y(PC[29]) );
  INVX12 U76 ( .A(n377), .Y(PC[30]) );
  AO21X4 U77 ( .A0(PCBrPredict[30]), .A1(n229), .B0(n261), .Y(n283) );
  INVX12 U78 ( .A(n50), .Y(PC[22]) );
  INVX12 U79 ( .A(n394), .Y(PC[24]) );
  INVX12 U80 ( .A(n54), .Y(PC[20]) );
  INVX12 U81 ( .A(n102), .Y(PC[10]) );
  INVX12 U82 ( .A(n106), .Y(PC[19]) );
  INVX12 U83 ( .A(n126), .Y(PC[16]) );
  INVX12 U84 ( .A(n184), .Y(PC[11]) );
  INVX12 U85 ( .A(n186), .Y(PC[14]) );
  INVX12 U86 ( .A(n188), .Y(PC[12]) );
  INVX12 U87 ( .A(n190), .Y(PC[18]) );
  INVX12 U88 ( .A(n192), .Y(PC[21]) );
  INVX12 U89 ( .A(n383), .Y(PC[17]) );
  INVX12 U90 ( .A(n196), .Y(PC[23]) );
  INVX12 U91 ( .A(n198), .Y(PC[9]) );
  OAI211X2 U92 ( .A0(n240), .A1(n303), .B0(n86), .C0(n87), .Y(n149) );
  INVX12 U93 ( .A(n200), .Y(PC[6]) );
  INVX12 U94 ( .A(n202), .Y(PC[7]) );
  INVX12 U95 ( .A(n204), .Y(PC[8]) );
  INVX12 U96 ( .A(n386), .Y(PC[13]) );
  INVX12 U97 ( .A(n208), .Y(PC[15]) );
  INVX1 U98 ( .A(n286), .Y(n279) );
  BUFX8 U99 ( .A(n279), .Y(n232) );
  NOR4X1 U100 ( .A(read_Instruction[5]), .B(read_Instruction[4]), .C(
        read_Instruction[31]), .D(read_Instruction[30]), .Y(n128) );
  INVX12 U101 ( .A(n210), .Y(PC[5]) );
  INVX12 U102 ( .A(n212), .Y(PC[4]) );
  INVX12 U103 ( .A(n214), .Y(n636) );
  INVX12 U104 ( .A(n216), .Y(PC[3]) );
  AND2X2 U106 ( .A(PCJumpJRorBranch[25]), .B(n231), .Y(n219) );
  NAND2X6 U107 ( .A(n222), .B(n20), .Y(n223) );
  AND2XL U108 ( .A(n285), .B(n319), .Y(n218) );
  CLKBUFX2 U109 ( .A(n19), .Y(n228) );
  CLKMX2X2 U110 ( .A(n518), .B(N25), .S0(n232), .Y(n220) );
  OAI2BB2X4 U111 ( .B0(n407), .B1(n123), .A0N(BranchTaken), .A1N(n123), .Y(
        next_BranchTaken) );
  NAND2X8 U112 ( .A(n223), .B(n242), .Y(n286) );
  AO22XL U113 ( .A0(Instruction[25]), .A1(n237), .B0(read_Instruction[25]), 
        .B1(n114), .Y(n182) );
  NAND3BXL U114 ( .AN(n234), .B(n263), .C(n262), .Y(n45) );
  NOR2X8 U115 ( .A(IF_ID_Write), .B(n286), .Y(n117) );
  AND4X4 U116 ( .A(n109), .B(n111), .C(n113), .D(next_BranchTaken), .Y(n121)
         );
  INVX1 U117 ( .A(PredictMiss), .Y(n257) );
  CLKINVX4 U118 ( .A(n125), .Y(n222) );
  CLKBUFX2 U119 ( .A(n19), .Y(n229) );
  CLKBUFX2 U120 ( .A(n278), .Y(n231) );
  OA21X4 U121 ( .A0(PredictMiss), .A1(IF_Flush), .B0(n242), .Y(n116) );
  NOR2XL U122 ( .A(n116), .B(n122), .Y(N109) );
  NOR2XL U123 ( .A(n112), .B(n116), .Y(N110) );
  NOR2XL U124 ( .A(n108), .B(n116), .Y(N114) );
  NOR2XL U125 ( .A(n111), .B(n116), .Y(N112) );
  NOR2XL U126 ( .A(n109), .B(n116), .Y(N113) );
  NOR2BXL U127 ( .AN(n113), .B(n116), .Y(N111) );
  CLKBUFX3 U128 ( .A(n224), .Y(n227) );
  NAND4XL U129 ( .A(n108), .B(n110), .C(n111), .D(n109), .Y(n256) );
  NOR2XL U130 ( .A(n112), .B(n113), .Y(n110) );
  CLKINVX1 U131 ( .A(stall), .Y(n242) );
  AOI22XL U132 ( .A0(Instruction[26]), .A1(n284), .B0(n117), .B1(
        read_Instruction[26]), .Y(n122) );
  AOI22X1 U133 ( .A0(n284), .A1(n584), .B0(n117), .B1(read_Instruction[27]), 
        .Y(n112) );
  AND2XL U134 ( .A(read_Instruction[14]), .B(n380), .Y(N175) );
  AND2XL U135 ( .A(read_Instruction[13]), .B(n380), .Y(N174) );
  AND2XL U136 ( .A(read_Instruction[12]), .B(n380), .Y(N173) );
  AND2XL U137 ( .A(read_Instruction[3]), .B(n380), .Y(N164) );
  AND2XL U138 ( .A(read_Instruction[4]), .B(n380), .Y(N165) );
  AND2XL U139 ( .A(read_Instruction[5]), .B(n380), .Y(N166) );
  AND2XL U140 ( .A(read_Instruction[6]), .B(n380), .Y(N167) );
  AND2XL U141 ( .A(read_Instruction[7]), .B(n380), .Y(N168) );
  AND2XL U142 ( .A(read_Instruction[8]), .B(n380), .Y(N169) );
  AND2XL U143 ( .A(read_Instruction[9]), .B(n380), .Y(N170) );
  AND2XL U144 ( .A(read_Instruction[10]), .B(n380), .Y(N171) );
  AND2XL U145 ( .A(read_Instruction[11]), .B(n380), .Y(N172) );
  INVXL U146 ( .A(read_Instruction[2]), .Y(n308) );
  AND2XL U147 ( .A(read_Instruction[1]), .B(n380), .Y(N162) );
  CLKAND2X3 U148 ( .A(read_Instruction[0]), .B(n380), .Y(N161) );
  INVXL U149 ( .A(read_Instruction[3]), .Y(n307) );
  INVXL U150 ( .A(read_Instruction[5]), .Y(n305) );
  AO22XL U151 ( .A0(read_Instruction[2]), .A1(n114), .B0(n418), .B1(n115), .Y(
        n159) );
  AO22XL U152 ( .A0(read_Instruction[4]), .A1(n114), .B0(n421), .B1(n237), .Y(
        n161) );
  AO22XL U153 ( .A0(read_Instruction[5]), .A1(n114), .B0(n437), .B1(n237), .Y(
        n162) );
  AO22XL U154 ( .A0(read_Instruction[0]), .A1(n114), .B0(Instruction[0]), .B1(
        n237), .Y(n157) );
  AO22XL U155 ( .A0(read_Instruction[1]), .A1(n114), .B0(Instruction[1]), .B1(
        n237), .Y(n158) );
  CLKMX2X2 U156 ( .A(n521), .B(N28), .S0(n232), .Y(n221) );
  INVXL U157 ( .A(read_Instruction[4]), .Y(n306) );
  INVXL U158 ( .A(read_Instruction[1]), .Y(n309) );
  INVX1 U159 ( .A(n105), .Y(n280) );
  INVX1 U160 ( .A(n104), .Y(n281) );
  AO22XL U161 ( .A0(Instruction[24]), .A1(n237), .B0(read_Instruction[24]), 
        .B1(n114), .Y(n181) );
  MX2XL U162 ( .A(n412), .B(N23), .S0(n232), .Y(n225) );
  MX2XL U163 ( .A(n415), .B(N24), .S0(n232), .Y(n226) );
  XNOR2XL U164 ( .A(n408), .B(PredictMiss), .Y(n119) );
  NAND2XL U165 ( .A(PredictMiss), .B(n287), .Y(n118) );
  INVX3 U166 ( .A(n241), .Y(n239) );
  INVX3 U167 ( .A(n241), .Y(n240) );
  CLKBUFX3 U168 ( .A(n243), .Y(n254) );
  CLKBUFX3 U169 ( .A(n243), .Y(n253) );
  CLKBUFX3 U170 ( .A(n245), .Y(n252) );
  CLKBUFX3 U171 ( .A(n244), .Y(n250) );
  CLKBUFX3 U172 ( .A(n244), .Y(n249) );
  CLKBUFX3 U173 ( .A(n245), .Y(n248) );
  CLKBUFX3 U174 ( .A(n244), .Y(n251) );
  CLKBUFX3 U175 ( .A(n243), .Y(n255) );
  INVX3 U177 ( .A(n235), .Y(n233) );
  CLKINVX1 U178 ( .A(n236), .Y(n234) );
  NAND2BX1 U179 ( .AN(n258), .B(n236), .Y(n259) );
  AOI2BB1X1 U180 ( .A0N(n263), .A1N(n257), .B0(IF_Flush), .Y(n258) );
  NOR2X1 U181 ( .A(n116), .B(n117), .Y(n115) );
  CLKINVX1 U182 ( .A(IF_Flush), .Y(n262) );
  CLKINVX1 U183 ( .A(n256), .Y(n263) );
  CLKBUFX3 U184 ( .A(n236), .Y(n235) );
  CLKBUFX3 U185 ( .A(n245), .Y(n247) );
  CLKBUFX3 U186 ( .A(n246), .Y(n245) );
  CLKBUFX3 U187 ( .A(n246), .Y(n243) );
  CLKBUFX3 U188 ( .A(n246), .Y(n244) );
  AOI2BB2X1 U189 ( .B0(PCBrPredict[29]), .B1(n229), .A0N(n240), .A1N(n264), 
        .Y(n265) );
  AOI2BB2X1 U190 ( .B0(PCJumpJRorBranch[29]), .B1(n231), .A0N(n235), .A1N(n397), .Y(n266) );
  CLKINVX1 U191 ( .A(n270), .Y(PCJumpEarly[27]) );
  CLKINVX1 U193 ( .A(n267), .Y(PCJumpEarly[28]) );
  CLKINVX1 U194 ( .A(n264), .Y(PCJumpEarly[29]) );
  CLKINVX1 U195 ( .A(n120), .Y(n287) );
  CLKINVX1 U196 ( .A(n285), .Y(n236) );
  NAND2BX1 U197 ( .AN(PCWrite), .B(n232), .Y(n285) );
  CLKBUFX3 U198 ( .A(rst), .Y(n246) );
  CLKINVX1 U199 ( .A(read_Instruction[6]), .Y(n304) );
  AOI22XL U200 ( .A0(PCBrPredict[8]), .A1(n228), .B0(n336), .B1(n233), .Y(n89)
         );
  NAND2X1 U201 ( .A(PCJumpJRorBranch[8]), .B(n231), .Y(n88) );
  CLKINVX1 U202 ( .A(read_Instruction[7]), .Y(n303) );
  AOI22XL U203 ( .A0(PCBrPredict[9]), .A1(n228), .B0(n335), .B1(n233), .Y(n87)
         );
  NAND2X1 U204 ( .A(PCJumpJRorBranch[9]), .B(n231), .Y(n86) );
  CLKINVX1 U205 ( .A(read_Instruction[8]), .Y(n302) );
  AOI22XL U206 ( .A0(PCBrPredict[10]), .A1(n228), .B0(n334), .B1(n233), .Y(n85) );
  NAND2X1 U207 ( .A(PCJumpJRorBranch[10]), .B(n231), .Y(n84) );
  CLKINVX1 U208 ( .A(read_Instruction[9]), .Y(n301) );
  AOI22XL U209 ( .A0(PCBrPredict[11]), .A1(n228), .B0(n333), .B1(n233), .Y(n83) );
  NAND2X1 U210 ( .A(PCJumpJRorBranch[11]), .B(n230), .Y(n82) );
  CLKINVX1 U211 ( .A(read_Instruction[10]), .Y(n300) );
  AOI22XL U212 ( .A0(PCBrPredict[12]), .A1(n228), .B0(n332), .B1(n233), .Y(n81) );
  NAND2X1 U213 ( .A(PCJumpJRorBranch[12]), .B(n278), .Y(n80) );
  OAI211X1 U214 ( .A0(n239), .A1(n299), .B0(n78), .C0(n79), .Y(n145) );
  CLKINVX1 U215 ( .A(read_Instruction[11]), .Y(n299) );
  AOI22XL U216 ( .A0(PCBrPredict[13]), .A1(n228), .B0(n385), .B1(n285), .Y(n79) );
  NAND2X1 U217 ( .A(PCJumpJRorBranch[13]), .B(n231), .Y(n78) );
  CLKINVX1 U218 ( .A(read_Instruction[12]), .Y(n298) );
  AOI22XL U219 ( .A0(PCBrPredict[14]), .A1(n228), .B0(n330), .B1(n233), .Y(n77) );
  NAND2X1 U220 ( .A(PCJumpJRorBranch[14]), .B(n278), .Y(n76) );
  OAI211X1 U221 ( .A0(n239), .A1(n297), .B0(n74), .C0(n75), .Y(n143) );
  CLKINVX1 U222 ( .A(read_Instruction[13]), .Y(n297) );
  AOI22XL U223 ( .A0(PCBrPredict[15]), .A1(n229), .B0(n329), .B1(n285), .Y(n75) );
  NAND2X1 U224 ( .A(PCJumpJRorBranch[15]), .B(n230), .Y(n74) );
  CLKINVX1 U225 ( .A(read_Instruction[14]), .Y(n296) );
  AOI22XL U226 ( .A0(PCBrPredict[16]), .A1(n19), .B0(n328), .B1(n233), .Y(n73)
         );
  NAND2X1 U227 ( .A(PCJumpJRorBranch[16]), .B(n230), .Y(n72) );
  CLKINVX1 U228 ( .A(read_Instruction[16]), .Y(n294) );
  AOI22XL U229 ( .A0(PCBrPredict[18]), .A1(n19), .B0(n326), .B1(n233), .Y(n69)
         );
  NAND2X1 U230 ( .A(PCJumpJRorBranch[18]), .B(n230), .Y(n68) );
  CLKINVX1 U231 ( .A(read_Instruction[17]), .Y(n293) );
  AOI22XL U232 ( .A0(PCBrPredict[19]), .A1(n19), .B0(n325), .B1(n233), .Y(n67)
         );
  NAND2X1 U233 ( .A(PCJumpJRorBranch[19]), .B(n230), .Y(n66) );
  CLKINVX1 U234 ( .A(read_Instruction[18]), .Y(n292) );
  AOI22XL U235 ( .A0(PCBrPredict[20]), .A1(n19), .B0(n324), .B1(n233), .Y(n65)
         );
  NAND2X1 U236 ( .A(PCJumpJRorBranch[20]), .B(n230), .Y(n64) );
  CLKINVX1 U237 ( .A(read_Instruction[19]), .Y(n291) );
  AOI22XL U238 ( .A0(PCBrPredict[21]), .A1(n19), .B0(n323), .B1(n233), .Y(n63)
         );
  NAND2X1 U239 ( .A(PCJumpJRorBranch[21]), .B(n230), .Y(n62) );
  CLKINVX1 U240 ( .A(read_Instruction[20]), .Y(n290) );
  AOI22XL U241 ( .A0(PCBrPredict[22]), .A1(n229), .B0(n322), .B1(n233), .Y(n61) );
  NAND2X1 U242 ( .A(PCJumpJRorBranch[22]), .B(n230), .Y(n60) );
  CLKINVX1 U243 ( .A(read_Instruction[21]), .Y(n289) );
  AOI22XL U244 ( .A0(PCBrPredict[23]), .A1(n229), .B0(n321), .B1(n234), .Y(n59) );
  NAND2X1 U245 ( .A(PCJumpJRorBranch[23]), .B(n230), .Y(n58) );
  CLKINVX1 U246 ( .A(read_Instruction[22]), .Y(n288) );
  AOI22XL U247 ( .A0(PCBrPredict[24]), .A1(n228), .B0(n387), .B1(n233), .Y(n57) );
  NAND2X1 U248 ( .A(PCJumpJRorBranch[24]), .B(n230), .Y(n56) );
  OAI211X1 U249 ( .A0(n240), .A1(n310), .B0(n100), .C0(n101), .Y(n156) );
  AOI22XL U250 ( .A0(PCBrPredict[2]), .A1(n228), .B0(n233), .B1(n636), .Y(n101) );
  NAND2X1 U251 ( .A(PCJumpJRorBranch[2]), .B(n231), .Y(n100) );
  OAI211X1 U252 ( .A0(n240), .A1(n309), .B0(n98), .C0(n99), .Y(n155) );
  AOI22XL U253 ( .A0(PCBrPredict[3]), .A1(n228), .B0(n341), .B1(n233), .Y(n99)
         );
  NAND2X1 U254 ( .A(PCJumpJRorBranch[3]), .B(n231), .Y(n98) );
  OAI211X1 U255 ( .A0(n240), .A1(n381), .B0(n96), .C0(n97), .Y(n154) );
  AOI22XL U256 ( .A0(PCBrPredict[4]), .A1(n228), .B0(PC[4]), .B1(n233), .Y(n97) );
  NAND2X1 U257 ( .A(PCJumpJRorBranch[4]), .B(n231), .Y(n96) );
  AOI22XL U258 ( .A0(PCBrPredict[7]), .A1(n228), .B0(n337), .B1(n233), .Y(n91)
         );
  NAND2X1 U259 ( .A(PCJumpJRorBranch[7]), .B(n278), .Y(n90) );
  CLKINVX1 U260 ( .A(read_Instruction[15]), .Y(n295) );
  AOI22XL U261 ( .A0(PCBrPredict[17]), .A1(n229), .B0(n382), .B1(n285), .Y(n71) );
  NAND2X1 U262 ( .A(PCJumpJRorBranch[17]), .B(n230), .Y(n70) );
  OAI211X1 U263 ( .A0(n307), .A1(n240), .B0(n94), .C0(n95), .Y(n153) );
  AOI22XL U264 ( .A0(PCBrPredict[5]), .A1(n228), .B0(n339), .B1(n233), .Y(n95)
         );
  NAND2X1 U265 ( .A(PCJumpJRorBranch[5]), .B(n231), .Y(n94) );
  AOI22XL U266 ( .A0(PCBrPredict[6]), .A1(n228), .B0(n338), .B1(n233), .Y(n93)
         );
  NAND2X1 U267 ( .A(PCJumpJRorBranch[6]), .B(n278), .Y(n92) );
  AOI2BB2X1 U268 ( .B0(PCBrPredict[26]), .B1(n229), .A0N(n240), .A1N(n273), 
        .Y(n274) );
  AOI2BB2X1 U269 ( .B0(PCJumpJRorBranch[26]), .B1(n230), .A0N(n235), .A1N(n400), .Y(n275) );
  AOI222XL U270 ( .A0(PC[0]), .A1(n233), .B0(PCJumpJRorBranch[0]), .B1(n230), 
        .C0(PCBrPredict[0]), .C1(n229), .Y(n105) );
  AOI222XL U271 ( .A0(PC[1]), .A1(n233), .B0(PCJumpJRorBranch[1]), .B1(n230), 
        .C0(PCBrPredict[1]), .C1(n229), .Y(n104) );
  AOI22X1 U272 ( .A0(n241), .A1(read_Instruction[23]), .B0(PCBrPredict[25]), 
        .B1(n229), .Y(n276) );
  AOI2BB2X1 U274 ( .B0(PCBrPredict[28]), .B1(n229), .A0N(n240), .A1N(n267), 
        .Y(n268) );
  AOI2BB2X1 U275 ( .B0(PCJumpJRorBranch[28]), .B1(n231), .A0N(n235), .A1N(n403), .Y(n269) );
  AOI2BB2X1 U276 ( .B0(PCBrPredict[27]), .B1(n229), .A0N(n240), .A1N(n270), 
        .Y(n271) );
  AO22X1 U279 ( .A0(read_Instruction[3]), .A1(n114), .B0(n488), .B1(n237), .Y(
        n160) );
  AO22X1 U280 ( .A0(read_Instruction[14]), .A1(n114), .B0(n459), .B1(n237), 
        .Y(n171) );
  AO22X1 U281 ( .A0(read_Instruction[13]), .A1(n114), .B0(n462), .B1(n237), 
        .Y(n170) );
  AO22X1 U282 ( .A0(read_Instruction[9]), .A1(n114), .B0(n430), .B1(n237), .Y(
        n166) );
  AO22X1 U283 ( .A0(read_Instruction[12]), .A1(n114), .B0(n456), .B1(n237), 
        .Y(n169) );
  AO22X1 U284 ( .A0(read_Instruction[8]), .A1(n114), .B0(n427), .B1(n237), .Y(
        n165) );
  AO22X1 U285 ( .A0(read_Instruction[11]), .A1(n114), .B0(n453), .B1(n237), 
        .Y(n168) );
  AO22X1 U286 ( .A0(read_Instruction[6]), .A1(n114), .B0(n424), .B1(n237), .Y(
        n163) );
  AO22X1 U287 ( .A0(read_Instruction[7]), .A1(n114), .B0(n441), .B1(n237), .Y(
        n164) );
  AO22X1 U288 ( .A0(read_Instruction[15]), .A1(n114), .B0(n444), .B1(n237), 
        .Y(n172) );
  AO22X1 U289 ( .A0(read_Instruction[10]), .A1(n114), .B0(Instruction[10]), 
        .B1(n237), .Y(n167) );
  AO22X1 U290 ( .A0(read_Instruction[16]), .A1(n114), .B0(Instruction[16]), 
        .B1(n237), .Y(n173) );
  AO22X1 U291 ( .A0(read_Instruction[17]), .A1(n114), .B0(Instruction[17]), 
        .B1(n237), .Y(n174) );
  AO22X1 U292 ( .A0(read_Instruction[18]), .A1(n114), .B0(Instruction[18]), 
        .B1(n237), .Y(n175) );
  AO22X1 U293 ( .A0(read_Instruction[19]), .A1(n114), .B0(Instruction[19]), 
        .B1(n237), .Y(n176) );
  AO22X1 U294 ( .A0(read_Instruction[20]), .A1(n114), .B0(Instruction[20]), 
        .B1(n237), .Y(n177) );
  AO22X1 U295 ( .A0(read_Instruction[21]), .A1(n114), .B0(Instruction[21]), 
        .B1(n237), .Y(n178) );
  AO22X1 U296 ( .A0(read_Instruction[22]), .A1(n114), .B0(Instruction[22]), 
        .B1(n237), .Y(n179) );
  AO22X1 U297 ( .A0(read_Instruction[23]), .A1(n114), .B0(Instruction[23]), 
        .B1(n237), .Y(n180) );
  AOI22X1 U298 ( .A0(Instruction[31]), .A1(n284), .B0(n117), .B1(
        read_Instruction[31]), .Y(n108) );
  AOI22X1 U299 ( .A0(Instruction[30]), .A1(n284), .B0(n117), .B1(
        read_Instruction[30]), .Y(n109) );
  AOI22X1 U300 ( .A0(Instruction[29]), .A1(n284), .B0(n117), .B1(
        read_Instruction[29]), .Y(n111) );
  AO22X1 U301 ( .A0(n284), .A1(Instruction[28]), .B0(n117), .B1(
        read_Instruction[28]), .Y(n113) );
  CLKINVX1 U302 ( .A(read_Instruction[0]), .Y(n310) );
  AND2X2 U303 ( .A(read_Instruction[2]), .B(n380), .Y(N163) );
  NOR3X1 U304 ( .A(Instruction[29]), .B(Instruction[31]), .C(Instruction[30]), 
        .Y(n124) );
  OAI22XL U305 ( .A0(n287), .A1(n8), .B0(n119), .B1(n120), .Y(N73) );
  OAI2BB2XL U306 ( .B0(n118), .B1(n8), .A0N(n118), .A1N(n407), .Y(N74) );
  InstructionFetch_DW01_add_0 add_71 ( .A({n313, n314, n315, n316, n317, n318, 
        n319, n387, n321, n322, n323, n324, n325, n326, n382, n328, n329, n330, 
        n385, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
        n13, n12}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), 
        .CI(1'b0), .SUM({N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, 
        N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, 
        N29, N28, N27, N26, N25, N24, N23}) );
  InstructionFetch_DW01_add_1 add_57_aco ( .A({PCJumpEarly[29:27], n384, n16, 
        n18, n17, n6, n5, n7, n4, n2, n9, n11, n10, n30, n27, n28, n29, n26, 
        n23, n24, n22, n25, n21, n15, n221, n14, n3, n220, n226, n225}), .B({
        n227, n227, n227, n227, n227, n227, n227, n224, n224, n227, n224, n227, 
        n227, n227, n224, N175, N174, N173, N172, N171, N170, N169, N168, N167, 
        N166, N165, N164, N163, N162, N161, 1'b0, 1'b0}), .CI(1'b0), .SUM(
        PCBrPredict) );
  TLATX1 \next_state_reg[0]  ( .G(n232), .D(N73), .Q(next_state[0]) );
  SDFFRX2 \PC_reg[31]  ( .D(n282), .SI(PC[30]), .SE(test_se), .CK(clk), .RN(
        n247), .Q(n313), .QN(n35) );
  SDFFRX2 \PC_reg[9]  ( .D(n149), .SI(PC[8]), .SE(test_se), .CK(clk), .RN(n248), .Q(n335), .QN(n198) );
  SDFFRX2 \PC_reg[3]  ( .D(n155), .SI(n636), .SE(test_se), .CK(clk), .RN(n249), 
        .Q(n341), .QN(n216) );
  SDFFRX2 \PC_reg[2]  ( .D(n156), .SI(n13), .SE(test_se), .CK(clk), .RN(n249), 
        .Q(n342), .QN(n214) );
  SDFFSXL \state_reg[0]  ( .D(next_state[0]), .SI(n51), .SE(test_se), .CK(clk), 
        .SN(n255), .Q(n376), .QN(n8) );
  SDFFRXL \Instruction_reg[1]  ( .D(n158), .SI(n374), .SE(test_se), .CK(clk), 
        .RN(n251), .Q(Instruction[1]), .QN(n375) );
  SDFFRXL \Instruction_reg[0]  ( .D(n157), .SI(n42), .SE(test_se), .CK(clk), 
        .RN(n252), .Q(Instruction[0]), .QN(n374) );
  SDFFRXL \Instruction_reg[10]  ( .D(n167), .SI(n364), .SE(test_se), .CK(clk), 
        .RN(n251), .Q(Instruction[10]), .QN(n373) );
  SDFFRXL \Instruction_reg[5]  ( .D(n162), .SI(n368), .SE(test_se), .CK(clk), 
        .RN(n251), .Q(n632), .QN(n372) );
  SDFFRXL \Instruction_reg[7]  ( .D(n164), .SI(n369), .SE(test_se), .CK(clk), 
        .RN(n251), .Q(n630), .QN(n371) );
  SDFFRXL \Instruction_reg[2]  ( .D(n159), .SI(n375), .SE(test_se), .CK(clk), 
        .RN(n251), .Q(n635), .QN(n370) );
  SDFFRXL \Instruction_reg[6]  ( .D(n163), .SI(n372), .SE(test_se), .CK(clk), 
        .RN(n251), .Q(n631), .QN(n369) );
  SDFFRXL \Instruction_reg[4]  ( .D(n161), .SI(n348), .SE(test_se), .CK(clk), 
        .RN(n251), .Q(n633), .QN(n368) );
  SDFFRXL \Instruction_reg[11]  ( .D(n168), .SI(n373), .SE(test_se), .CK(clk), 
        .RN(n251), .Q(n627), .QN(n367) );
  SDFFRXL \Instruction_reg[8]  ( .D(n165), .SI(n371), .SE(test_se), .CK(clk), 
        .RN(n251), .Q(n629), .QN(n366) );
  SDFFRXL \Instruction_reg[12]  ( .D(n169), .SI(n367), .SE(test_se), .CK(clk), 
        .RN(n250), .Q(n626), .QN(n365) );
  SDFFRXL \Instruction_reg[9]  ( .D(n166), .SI(n366), .SE(test_se), .CK(clk), 
        .RN(n251), .Q(n628), .QN(n364) );
  SDFFSXL \state_reg[1]  ( .D(next_state[1]), .SI(n376), .SE(test_se), .CK(clk), .SN(n255), .Q(\state[1] ), .QN(test_so) );
  SDFFRXL \PCadd4_reg[1]  ( .D(n226), .SI(n361), .SE(test_se), .CK(clk), .RN(
        n254), .Q(n615), .QN(n362) );
  SDFFRXL \PCadd4_reg[0]  ( .D(n225), .SI(PC[31]), .SE(test_se), .CK(clk), 
        .RN(n255), .Q(n616), .QN(n361) );
  SDFFRXL \Instruction_reg[23]  ( .D(n180), .SI(n359), .SE(test_se), .CK(clk), 
        .RN(n250), .Q(Instruction[23]), .QN(n360) );
  SDFFRXL \Instruction_reg[22]  ( .D(n179), .SI(n358), .SE(test_se), .CK(clk), 
        .RN(n250), .Q(Instruction[22]), .QN(n359) );
  SDFFRXL \Instruction_reg[21]  ( .D(n178), .SI(n357), .SE(test_se), .CK(clk), 
        .RN(n250), .Q(Instruction[21]), .QN(n358) );
  SDFFRXL \Instruction_reg[20]  ( .D(n177), .SI(n356), .SE(test_se), .CK(clk), 
        .RN(n250), .Q(Instruction[20]), .QN(n357) );
  SDFFRXL \Instruction_reg[19]  ( .D(n176), .SI(n355), .SE(test_se), .CK(clk), 
        .RN(n250), .Q(Instruction[19]), .QN(n356) );
  SDFFRXL \Instruction_reg[18]  ( .D(n175), .SI(n354), .SE(test_se), .CK(clk), 
        .RN(n250), .Q(Instruction[18]), .QN(n355) );
  SDFFRXL \Instruction_reg[17]  ( .D(n174), .SI(n353), .SE(test_se), .CK(clk), 
        .RN(n250), .Q(Instruction[17]), .QN(n354) );
  SDFFRXL \Instruction_reg[16]  ( .D(n173), .SI(n49), .SE(test_se), .CK(clk), 
        .RN(n250), .Q(Instruction[16]), .QN(n353) );
  SDFFRXL \Instruction_reg[25]  ( .D(n182), .SI(n351), .SE(test_se), .CK(clk), 
        .RN(n249), .Q(Instruction[25]), .QN(n352) );
  SDFFRXL \Instruction_reg[24]  ( .D(n181), .SI(n360), .SE(test_se), .CK(clk), 
        .RN(n249), .Q(Instruction[24]), .QN(n351) );
  SDFFRXL \Instruction_reg[13]  ( .D(n170), .SI(n365), .SE(test_se), .CK(clk), 
        .RN(n250), .Q(n625), .QN(n350) );
  SDFFRXL \Instruction_reg[14]  ( .D(n171), .SI(n350), .SE(test_se), .CK(clk), 
        .RN(n250), .Q(n624), .QN(n349) );
  SDFFRXL \Instruction_reg[3]  ( .D(n160), .SI(n370), .SE(test_se), .CK(clk), 
        .RN(n251), .Q(n634), .QN(n348) );
  SDFFRXL \PCadd4_reg[27]  ( .D(n16), .SI(n346), .SE(test_se), .CK(clk), .RN(
        n252), .Q(n589), .QN(n347) );
  SDFFRXL \PCadd4_reg[26]  ( .D(n18), .SI(n345), .SE(test_se), .CK(clk), .RN(
        n252), .Q(n590), .QN(n346) );
  SDFFRXL \PCadd4_reg[25]  ( .D(n17), .SI(n344), .SE(test_se), .CK(clk), .RN(
        n252), .Q(n591), .QN(n345) );
  SDFFRXL \PCadd4_reg[24]  ( .D(n6), .SI(n343), .SE(test_se), .CK(clk), .RN(
        n253), .Q(n592), .QN(n344) );
  SDFFRXL \PCadd4_reg[23]  ( .D(n5), .SI(n312), .SE(test_se), .CK(clk), .RN(
        n253), .Q(n593), .QN(n343) );
  SDFFRXL \PCadd4_reg[22]  ( .D(n7), .SI(n311), .SE(test_se), .CK(clk), .RN(
        n253), .Q(n594), .QN(n312) );
  SDFFRXL \PCadd4_reg[21]  ( .D(n4), .SI(n217), .SE(test_se), .CK(clk), .RN(
        n253), .Q(n595), .QN(n311) );
  SDFFRXL \PCadd4_reg[20]  ( .D(n2), .SI(n215), .SE(test_se), .CK(clk), .RN(
        n253), .Q(n596), .QN(n217) );
  SDFFRXL \PCadd4_reg[19]  ( .D(n9), .SI(n213), .SE(test_se), .CK(clk), .RN(
        n253), .Q(n597), .QN(n215) );
  SDFFRXL \PCadd4_reg[18]  ( .D(n11), .SI(n211), .SE(test_se), .CK(clk), .RN(
        n253), .Q(n598), .QN(n213) );
  SDFFRXL \PCadd4_reg[17]  ( .D(n10), .SI(n209), .SE(test_se), .CK(clk), .RN(
        n253), .Q(n599), .QN(n211) );
  SDFFRXL \PCadd4_reg[16]  ( .D(n30), .SI(n207), .SE(test_se), .CK(clk), .RN(
        n253), .Q(n600), .QN(n209) );
  SDFFRXL \PCadd4_reg[15]  ( .D(n27), .SI(n205), .SE(test_se), .CK(clk), .RN(
        n253), .Q(n601), .QN(n207) );
  SDFFRXL \PCadd4_reg[14]  ( .D(n28), .SI(n203), .SE(test_se), .CK(clk), .RN(
        n253), .Q(n602), .QN(n205) );
  SDFFRXL \PCadd4_reg[13]  ( .D(n29), .SI(n201), .SE(test_se), .CK(clk), .RN(
        n253), .Q(n603), .QN(n203) );
  SDFFRXL \PCadd4_reg[12]  ( .D(n26), .SI(n199), .SE(test_se), .CK(clk), .RN(
        n254), .Q(n604), .QN(n201) );
  SDFFRXL \PCadd4_reg[11]  ( .D(n23), .SI(n197), .SE(test_se), .CK(clk), .RN(
        n254), .Q(n605), .QN(n199) );
  SDFFRXL \PCadd4_reg[10]  ( .D(n24), .SI(n195), .SE(test_se), .CK(clk), .RN(
        n254), .Q(n606), .QN(n197) );
  SDFFRXL \PCadd4_reg[9]  ( .D(n22), .SI(n193), .SE(test_se), .CK(clk), .RN(
        n254), .Q(n607), .QN(n195) );
  SDFFRXL \PCadd4_reg[8]  ( .D(n25), .SI(n191), .SE(test_se), .CK(clk), .RN(
        n254), .Q(n608), .QN(n193) );
  SDFFRXL \PCadd4_reg[7]  ( .D(n21), .SI(n189), .SE(test_se), .CK(clk), .RN(
        n254), .Q(n609), .QN(n191) );
  SDFFRXL \PCadd4_reg[6]  ( .D(n15), .SI(n187), .SE(test_se), .CK(clk), .RN(
        n254), .Q(n610), .QN(n189) );
  SDFFRXL \PCadd4_reg[5]  ( .D(n221), .SI(n185), .SE(test_se), .CK(clk), .RN(
        n254), .Q(n611), .QN(n187) );
  SDFFRXL \PCadd4_reg[4]  ( .D(n14), .SI(n183), .SE(test_se), .CK(clk), .RN(
        n254), .Q(n612), .QN(n185) );
  SDFFRXL \PCadd4_reg[3]  ( .D(n3), .SI(n107), .SE(test_se), .CK(clk), .RN(
        n254), .Q(n613), .QN(n183) );
  SDFFRXL \PCadd4_reg[2]  ( .D(n220), .SI(n362), .SE(test_se), .CK(clk), .RN(
        n254), .Q(n614), .QN(n107) );
  SDFFRXL \PCadd4_reg[28]  ( .D(n384), .SI(n347), .SE(test_se), .CK(clk), .RN(
        n252), .Q(n588), .QN(n103) );
  SDFFRXL \PCadd4_reg[29]  ( .D(PCJumpEarly[27]), .SI(n103), .SE(test_se), 
        .CK(clk), .RN(n252), .Q(n587), .QN(n55) );
  SDFFRXL \PCadd4_reg[30]  ( .D(PCJumpEarly[28]), .SI(n55), .SE(test_se), .CK(
        clk), .RN(n252), .Q(n586), .QN(n53) );
  SDFFRXL \PCadd4_reg[31]  ( .D(PCJumpEarly[29]), .SI(n53), .SE(test_se), .CK(
        clk), .RN(n252), .Q(n585), .QN(n51) );
  SDFFRXL \Instruction_reg[15]  ( .D(n172), .SI(n349), .SE(test_se), .CK(clk), 
        .RN(n250), .Q(n623), .QN(n49) );
  SDFFRXL \Instruction_reg[29]  ( .D(N112), .SI(n36), .SE(test_se), .CK(clk), 
        .RN(n247), .Q(n619), .QN(n47) );
  SDFFRXL \Instruction_reg[30]  ( .D(N113), .SI(n47), .SE(test_se), .CK(clk), 
        .RN(n247), .Q(n618), .QN(n44) );
  SDFFRXL \PC_reg[30]  ( .D(n283), .SI(PC[29]), .SE(test_se), .CK(clk), .RN(
        n247), .Q(n314), .QN(n48) );
  SDFFRXL \PC_reg[0]  ( .D(n280), .SI(n34), .SE(test_se), .CK(clk), .RN(n249), 
        .Q(n12), .QN(n31) );
  SDFFRXL \PC_reg[1]  ( .D(n281), .SI(n12), .SE(test_se), .CK(clk), .RN(n249), 
        .Q(n13), .QN(n32) );
  SDFFRXL BranchTaken_reg ( .D(next_BranchTaken), .SI(test_si), .SE(test_se), 
        .CK(clk), .RN(n249), .Q(BranchTaken), .QN(n42) );
  SDFFRXL \Instruction_reg[27]  ( .D(N110), .SI(n38), .SE(test_se), .CK(clk), 
        .RN(n247), .Q(n621), .QN(n40) );
  SDFFRXL \Instruction_reg[26]  ( .D(N109), .SI(n352), .SE(test_se), .CK(clk), 
        .RN(n249), .Q(n622), .QN(n38) );
  SDFFRXL \Instruction_reg[28]  ( .D(N111), .SI(n40), .SE(test_se), .CK(clk), 
        .RN(n247), .Q(n620), .QN(n36) );
  SDFFRXL \Instruction_reg[31]  ( .D(N114), .SI(n44), .SE(test_se), .CK(clk), 
        .RN(n251), .Q(n617), .QN(n34) );
  SDFFRXL \PC_reg[27]  ( .D(n131), .SI(PC[26]), .SE(test_se), .CK(clk), .RN(
        n252), .Q(n317), .QN(n39) );
  SDFFRXL \PC_reg[28]  ( .D(n130), .SI(PC[27]), .SE(test_se), .CK(clk), .RN(
        n252), .Q(n316), .QN(n43) );
  SDFFRXL \PC_reg[26]  ( .D(n132), .SI(PC[25]), .SE(test_se), .CK(clk), .RN(
        n252), .Q(n318), .QN(n41) );
  SDFFRXL \PC_reg[29]  ( .D(n129), .SI(PC[28]), .SE(test_se), .CK(clk), .RN(
        n252), .Q(n315), .QN(n46) );
  SDFFRXL \PC_reg[25]  ( .D(n133), .SI(PC[24]), .SE(test_se), .CK(clk), .RN(
        n247), .Q(n319), .QN(n37) );
  SDFFRXL \PC_reg[23]  ( .D(n135), .SI(PC[22]), .SE(test_se), .CK(clk), .RN(
        n247), .Q(n321), .QN(n196) );
  SDFFRXL \PC_reg[22]  ( .D(n136), .SI(PC[21]), .SE(test_se), .CK(clk), .RN(
        n247), .Q(n322), .QN(n50) );
  SDFFRXL \PC_reg[21]  ( .D(n137), .SI(PC[20]), .SE(test_se), .CK(clk), .RN(
        n247), .Q(n323), .QN(n192) );
  SDFFRXL \PC_reg[20]  ( .D(n138), .SI(PC[19]), .SE(test_se), .CK(clk), .RN(
        n247), .Q(n324), .QN(n54) );
  SDFFRXL \PC_reg[19]  ( .D(n139), .SI(PC[18]), .SE(test_se), .CK(clk), .RN(
        n248), .Q(n325), .QN(n106) );
  SDFFRXL \PC_reg[18]  ( .D(n140), .SI(PC[17]), .SE(test_se), .CK(clk), .RN(
        n248), .Q(n326), .QN(n190) );
  SDFFRXL \PC_reg[16]  ( .D(n142), .SI(PC[15]), .SE(test_se), .CK(clk), .RN(
        n248), .Q(n328), .QN(n126) );
  SDFFRXL \PC_reg[15]  ( .D(n143), .SI(PC[14]), .SE(test_se), .CK(clk), .RN(
        n248), .Q(n329), .QN(n208) );
  SDFFRXL \PC_reg[14]  ( .D(n144), .SI(PC[13]), .SE(test_se), .CK(clk), .RN(
        n248), .Q(n330), .QN(n186) );
  SDFFRXL \PC_reg[12]  ( .D(n146), .SI(PC[11]), .SE(test_se), .CK(clk), .RN(
        n248), .Q(n332), .QN(n188) );
  SDFFRXL \PC_reg[11]  ( .D(n147), .SI(PC[10]), .SE(test_se), .CK(clk), .RN(
        n248), .Q(n333), .QN(n184) );
  SDFFRXL \PC_reg[10]  ( .D(n148), .SI(PC[9]), .SE(test_se), .CK(clk), .RN(
        n248), .Q(n334), .QN(n102) );
  SDFFRXL \PC_reg[8]  ( .D(n150), .SI(PC[7]), .SE(test_se), .CK(clk), .RN(n248), .Q(n336), .QN(n204) );
  SDFFRXL \PC_reg[7]  ( .D(n151), .SI(PC[6]), .SE(test_se), .CK(clk), .RN(n249), .Q(n337), .QN(n202) );
  SDFFRXL \PC_reg[6]  ( .D(n152), .SI(PC[5]), .SE(test_se), .CK(clk), .RN(n249), .Q(n338), .QN(n200) );
  SDFFRXL \PC_reg[5]  ( .D(n153), .SI(n340), .SE(test_se), .CK(clk), .RN(n249), 
        .Q(n339), .QN(n210) );
  SDFFRXL \PC_reg[4]  ( .D(n154), .SI(PC[3]), .SE(test_se), .CK(clk), .RN(n249), .Q(n340), .QN(n212) );
  SDFFRX4 \PC_reg[24]  ( .D(n134), .SI(PC[23]), .SE(test_se), .CK(clk), .RN(
        n247), .Q(n387) );
  SDFFRHQX8 \PC_reg[13]  ( .D(n145), .SI(PC[12]), .SE(test_se), .CK(clk), .RN(
        n248), .Q(n385) );
  SDFFRHQX8 \PC_reg[17]  ( .D(n141), .SI(PC[16]), .SE(test_se), .CK(clk), .RN(
        n248), .Q(n382) );
  CLKBUFX2 U1 ( .A(n48), .Y(n377) );
  CLKBUFX2 U2 ( .A(n218), .Y(n378) );
  CLKBUFX2 U6 ( .A(n39), .Y(n379) );
  CLKBUFX20 U28 ( .A(N13), .Y(n380) );
  INVXL U60 ( .A(read_Instruction[2]), .Y(n381) );
  CLKINVX20 U66 ( .A(n382), .Y(n383) );
  CLKMX2X6 U105 ( .A(N51), .B(n497), .S0(n286), .Y(n384) );
  CLKINVX20 U176 ( .A(n384), .Y(n273) );
  CLKINVX20 U192 ( .A(n385), .Y(n386) );
  AOI22X4 U273 ( .A0(PCJumpJRorBranch[27]), .A1(n230), .B0(n390), .B1(n389), 
        .Y(n272) );
  CLKINVX20 U277 ( .A(n379), .Y(n389) );
  CLKINVX20 U278 ( .A(n235), .Y(n390) );
  OAI2BB2X4 U307 ( .B0(n35), .B1(n235), .A0N(PCJumpJRorBranch[31]), .A1N(n231), 
        .Y(n260) );
  OAI2BB2X4 U308 ( .B0(n377), .B1(n235), .A0N(PCJumpJRorBranch[30]), .A1N(n231), .Y(n261) );
  OR2X8 U309 ( .A(n237), .B(n116), .Y(n391) );
  CLKINVX20 U310 ( .A(n391), .Y(n114) );
  CLKINVX20 U311 ( .A(n378), .Y(n392) );
  OR2X8 U312 ( .A(n393), .B(n219), .Y(n133) );
  NAND2X8 U313 ( .A(n392), .B(n276), .Y(n393) );
  CLKINVX20 U314 ( .A(n387), .Y(n394) );
  INVXL U315 ( .A(n46), .Y(n395) );
  INVXL U316 ( .A(n395), .Y(n396) );
  INVXL U317 ( .A(n395), .Y(n397) );
  INVXL U318 ( .A(n41), .Y(n398) );
  INVXL U319 ( .A(n398), .Y(n399) );
  INVXL U320 ( .A(n398), .Y(n400) );
  INVXL U321 ( .A(n43), .Y(n401) );
  INVXL U322 ( .A(n401), .Y(n402) );
  INVXL U323 ( .A(n401), .Y(n403) );
  INVXL U324 ( .A(n39), .Y(n404) );
  INVXL U325 ( .A(n404), .Y(n405) );
  INVXL U326 ( .A(\state[1] ), .Y(n406) );
  INVXL U327 ( .A(n406), .Y(n407) );
  INVXL U328 ( .A(n406), .Y(n408) );
  CLKBUFX2 U329 ( .A(n484), .Y(PCadd4[29]) );
  INVXL U330 ( .A(n616), .Y(n410) );
  INVXL U331 ( .A(n410), .Y(PCadd4[0]) );
  INVXL U332 ( .A(n410), .Y(n412) );
  INVXL U333 ( .A(n615), .Y(n413) );
  INVXL U334 ( .A(n413), .Y(PCadd4[1]) );
  INVXL U335 ( .A(n413), .Y(n415) );
  INVXL U336 ( .A(n635), .Y(n416) );
  INVXL U337 ( .A(n416), .Y(Instruction[2]) );
  INVXL U338 ( .A(n416), .Y(n418) );
  INVXL U339 ( .A(n633), .Y(n419) );
  INVXL U340 ( .A(n419), .Y(Instruction[4]) );
  INVXL U341 ( .A(n419), .Y(n421) );
  INVXL U342 ( .A(n631), .Y(n422) );
  INVXL U343 ( .A(n422), .Y(Instruction[6]) );
  INVXL U344 ( .A(n422), .Y(n424) );
  INVXL U345 ( .A(n629), .Y(n425) );
  INVXL U346 ( .A(n425), .Y(Instruction[8]) );
  INVXL U347 ( .A(n425), .Y(n427) );
  INVXL U348 ( .A(n628), .Y(n428) );
  INVXL U349 ( .A(n428), .Y(Instruction[9]) );
  INVXL U350 ( .A(n428), .Y(n430) );
  CLKBUFX2 U351 ( .A(n499), .Y(PCadd4[27]) );
  CLKBUFX2 U352 ( .A(n491), .Y(PCadd4[3]) );
  CLKBUFX2 U353 ( .A(n493), .Y(PCadd4[31]) );
  CLKBUFX2 U354 ( .A(n496), .Y(PCadd4[28]) );
  INVXL U355 ( .A(n632), .Y(n435) );
  INVXL U356 ( .A(n435), .Y(Instruction[5]) );
  INVXL U357 ( .A(n435), .Y(n437) );
  CLKBUFX2 U358 ( .A(n487), .Y(Instruction[3]) );
  INVXL U359 ( .A(n630), .Y(n439) );
  INVXL U360 ( .A(n439), .Y(Instruction[7]) );
  INVXL U361 ( .A(n439), .Y(n441) );
  INVXL U362 ( .A(n623), .Y(n442) );
  INVXL U363 ( .A(n442), .Y(Instruction[15]) );
  INVXL U364 ( .A(n442), .Y(n444) );
  CLKBUFX2 U365 ( .A(n502), .Y(PCadd4[30]) );
  CLKBUFX2 U366 ( .A(n505), .Y(PCadd4[8]) );
  CLKBUFX2 U367 ( .A(n508), .Y(PCadd4[22]) );
  CLKBUFX2 U368 ( .A(n511), .Y(PCadd4[26]) );
  INVX12 U369 ( .A(n214), .Y(PC[2]) );
  CLKBUFX2 U370 ( .A(n517), .Y(PCadd4[2]) );
  INVXL U371 ( .A(n627), .Y(n451) );
  INVXL U372 ( .A(n451), .Y(Instruction[11]) );
  INVXL U373 ( .A(n451), .Y(n453) );
  INVXL U374 ( .A(n626), .Y(n454) );
  INVXL U375 ( .A(n454), .Y(Instruction[12]) );
  INVXL U376 ( .A(n454), .Y(n456) );
  INVXL U377 ( .A(n624), .Y(n457) );
  INVXL U378 ( .A(n457), .Y(Instruction[14]) );
  INVXL U379 ( .A(n457), .Y(n459) );
  INVXL U380 ( .A(n625), .Y(n460) );
  INVXL U381 ( .A(n460), .Y(Instruction[13]) );
  INVXL U382 ( .A(n460), .Y(n462) );
  CLKBUFX2 U383 ( .A(n514), .Y(PCadd4[21]) );
  CLKBUFX2 U384 ( .A(n520), .Y(PCadd4[5]) );
  CLKBUFX2 U385 ( .A(n523), .Y(PCadd4[9]) );
  CLKBUFX2 U386 ( .A(n526), .Y(PCadd4[11]) );
  CLKBUFX2 U387 ( .A(n529), .Y(PCadd4[13]) );
  CLKBUFX2 U388 ( .A(n532), .Y(PCadd4[17]) );
  CLKBUFX2 U389 ( .A(n535), .Y(PCadd4[4]) );
  CLKBUFX2 U390 ( .A(n544), .Y(PCadd4[6]) );
  CLKBUFX2 U391 ( .A(n547), .Y(PCadd4[12]) );
  CLKBUFX2 U392 ( .A(n550), .Y(PCadd4[14]) );
  CLKBUFX2 U393 ( .A(n553), .Y(PCadd4[18]) );
  CLKBUFX2 U394 ( .A(n538), .Y(PCadd4[23]) );
  CLKBUFX2 U395 ( .A(n541), .Y(PCadd4[24]) );
  CLKBUFX2 U396 ( .A(n556), .Y(PCadd4[16]) );
  CLKBUFX2 U397 ( .A(n559), .Y(PCadd4[19]) );
  CLKBUFX2 U398 ( .A(n562), .Y(PCadd4[25]) );
  CLKBUFX2 U399 ( .A(n565), .Y(PCadd4[10]) );
  CLKBUFX2 U400 ( .A(n568), .Y(PCadd4[20]) );
  CLKBUFX2 U401 ( .A(n572), .Y(PCadd4[7]) );
  CLKBUFX2 U402 ( .A(n574), .Y(PCadd4[15]) );
  INVXL U403 ( .A(n587), .Y(n483) );
  INVXL U404 ( .A(n483), .Y(n484) );
  INVXL U405 ( .A(n483), .Y(n485) );
  INVXL U406 ( .A(n634), .Y(n486) );
  INVXL U407 ( .A(n486), .Y(n487) );
  INVXL U408 ( .A(n486), .Y(n488) );
  INVXL U409 ( .A(n613), .Y(n489) );
  INVXL U410 ( .A(n489), .Y(n490) );
  INVXL U411 ( .A(n489), .Y(n491) );
  INVXL U412 ( .A(n585), .Y(n492) );
  INVXL U413 ( .A(n492), .Y(n493) );
  INVXL U414 ( .A(n492), .Y(n494) );
  INVXL U415 ( .A(n588), .Y(n495) );
  INVXL U416 ( .A(n495), .Y(n496) );
  INVXL U417 ( .A(n495), .Y(n497) );
  INVXL U418 ( .A(n589), .Y(n498) );
  INVXL U419 ( .A(n498), .Y(n499) );
  INVXL U420 ( .A(n498), .Y(n500) );
  INVXL U421 ( .A(n586), .Y(n501) );
  INVXL U422 ( .A(n501), .Y(n502) );
  INVXL U423 ( .A(n501), .Y(n503) );
  INVXL U424 ( .A(n608), .Y(n504) );
  INVXL U425 ( .A(n504), .Y(n505) );
  INVXL U426 ( .A(n504), .Y(n506) );
  INVXL U427 ( .A(n594), .Y(n507) );
  INVXL U428 ( .A(n507), .Y(n508) );
  INVXL U429 ( .A(n507), .Y(n509) );
  INVXL U430 ( .A(n590), .Y(n510) );
  INVXL U431 ( .A(n510), .Y(n511) );
  INVXL U432 ( .A(n510), .Y(n512) );
  INVXL U433 ( .A(n595), .Y(n513) );
  INVXL U434 ( .A(n513), .Y(n514) );
  INVXL U435 ( .A(n513), .Y(n515) );
  INVXL U436 ( .A(n614), .Y(n516) );
  INVXL U437 ( .A(n516), .Y(n517) );
  INVXL U438 ( .A(n516), .Y(n518) );
  INVXL U439 ( .A(n611), .Y(n519) );
  INVXL U440 ( .A(n519), .Y(n520) );
  INVXL U441 ( .A(n519), .Y(n521) );
  INVXL U442 ( .A(n607), .Y(n522) );
  INVXL U443 ( .A(n522), .Y(n523) );
  INVXL U444 ( .A(n522), .Y(n524) );
  INVXL U445 ( .A(n605), .Y(n525) );
  INVXL U446 ( .A(n525), .Y(n526) );
  INVXL U447 ( .A(n525), .Y(n527) );
  INVXL U448 ( .A(n603), .Y(n528) );
  INVXL U449 ( .A(n528), .Y(n529) );
  INVXL U450 ( .A(n528), .Y(n530) );
  INVXL U451 ( .A(n599), .Y(n531) );
  INVXL U452 ( .A(n531), .Y(n532) );
  INVXL U453 ( .A(n531), .Y(n533) );
  INVXL U454 ( .A(n612), .Y(n534) );
  INVXL U455 ( .A(n534), .Y(n535) );
  INVXL U456 ( .A(n534), .Y(n536) );
  INVXL U457 ( .A(n593), .Y(n537) );
  INVXL U458 ( .A(n537), .Y(n538) );
  INVXL U459 ( .A(n537), .Y(n539) );
  INVXL U460 ( .A(n592), .Y(n540) );
  INVXL U461 ( .A(n540), .Y(n541) );
  INVXL U462 ( .A(n540), .Y(n542) );
  INVXL U463 ( .A(n610), .Y(n543) );
  INVXL U464 ( .A(n543), .Y(n544) );
  INVXL U465 ( .A(n543), .Y(n545) );
  INVXL U466 ( .A(n604), .Y(n546) );
  INVXL U467 ( .A(n546), .Y(n547) );
  INVXL U468 ( .A(n546), .Y(n548) );
  INVXL U469 ( .A(n602), .Y(n549) );
  INVXL U470 ( .A(n549), .Y(n550) );
  INVXL U471 ( .A(n549), .Y(n551) );
  INVXL U472 ( .A(n598), .Y(n552) );
  INVXL U473 ( .A(n552), .Y(n553) );
  INVXL U474 ( .A(n552), .Y(n554) );
  INVXL U475 ( .A(n600), .Y(n555) );
  INVXL U476 ( .A(n555), .Y(n556) );
  INVXL U477 ( .A(n555), .Y(n557) );
  INVXL U478 ( .A(n597), .Y(n558) );
  INVXL U479 ( .A(n558), .Y(n559) );
  INVXL U480 ( .A(n558), .Y(n560) );
  INVXL U481 ( .A(n591), .Y(n561) );
  INVXL U482 ( .A(n561), .Y(n562) );
  INVXL U483 ( .A(n561), .Y(n563) );
  INVXL U484 ( .A(n606), .Y(n564) );
  INVXL U485 ( .A(n564), .Y(n565) );
  INVXL U486 ( .A(n564), .Y(n566) );
  INVXL U487 ( .A(n596), .Y(n567) );
  INVXL U488 ( .A(n567), .Y(n568) );
  INVXL U489 ( .A(n567), .Y(n569) );
  INVXL U490 ( .A(n609), .Y(n570) );
  INVXL U491 ( .A(n570), .Y(n571) );
  INVXL U492 ( .A(n570), .Y(n572) );
  INVXL U493 ( .A(n601), .Y(n573) );
  INVXL U494 ( .A(n573), .Y(n574) );
  INVXL U495 ( .A(n573), .Y(n575) );
  CLKBUFX2 U496 ( .A(n619), .Y(Instruction[29]) );
  CLKBUFX2 U497 ( .A(n618), .Y(Instruction[30]) );
  CLKBUFX2 U498 ( .A(n617), .Y(Instruction[31]) );
  CLKBUFX2 U499 ( .A(n620), .Y(Instruction[28]) );
  CLKBUFX2 U500 ( .A(n622), .Y(Instruction[26]) );
  CLKBUFX2 U501 ( .A(n583), .Y(Instruction[27]) );
  INVXL U502 ( .A(n621), .Y(n582) );
  INVXL U503 ( .A(n582), .Y(n583) );
  INVXL U504 ( .A(n582), .Y(n584) );
endmodule


module MIPS_Pipeline ( clk, rst, ICACHE_addr, ICACHE_rdata, ICACHE_ren, 
        ICACHE_wen, ICACHE_wdata, ICACHE_stall, DCACHE_addr, DCACHE_rdata, 
        DCACHE_ren, DCACHE_wen, DCACHE_wdata, DCACHE_stall, test_si, test_so, 
        test_se );
  output [31:0] ICACHE_addr;
  input [31:0] ICACHE_rdata;
  output [31:0] ICACHE_wdata;
  output [31:0] DCACHE_addr;
  input [31:0] DCACHE_rdata;
  output [31:0] DCACHE_wdata;
  input clk, rst, ICACHE_stall, DCACHE_stall, test_si, test_se;
  output ICACHE_ren, ICACHE_wen, DCACHE_ren, DCACHE_wen, test_so;
  wire   needStall, IF_Flush, PredictMiss, BranchTaken, PCBuffer_valid, Jump,
         Branch, \ALUOp[0] , ALUSrc, N182, N199, N202, n54, n55, n56, n57, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n237, n238, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         SYNOPSYS_UNCONNECTED__0, n3, n4, n5, n6;
  wire   [2:0] EX_MEM_MEMControl;
  wire   [31:0] PCJump_JRChecked;
  wire   [31:0] PCadd4;
  wire   [31:0] Instruction;
  wire   [31:0] PCbranched;
  wire   [4:0] MEM_WB_RegisterRd;
  wire   [1:0] ID_EX_WBControl;
  wire   [2:0] ID_EX_MEMControl;
  wire   [6:0] ID_EX_EXControl;
  wire   [31:0] ReadData1;
  wire   [31:0] ReadData2;
  wire   [31:0] next_ReadData1;
  wire   [31:0] Immediate_SE;
  wire   [4:0] ID_EX_RegisterRd;
  wire   [4:0] ID_EX_RegisterRs;
  wire   [4:0] ID_EX_RegisterRt;
  wire   [1:0] MEM_WB_WBControl;
  wire   [31:0] next_ALUresult;
  wire   [1:0] BrForwardA;
  wire   [1:0] BrForwardB;
  wire   [1:0] EX_MEM_WBControl;
  wire   [4:0] EX_MEM_RegisterRd;
  wire   [1:0] ForwardA;
  wire   [1:0] ForwardB;
  wire   [31:0] MemoryData;
  wire   [31:0] Buf_ALUresult;
  assign ICACHE_wdata[0] = 1'b0;
  assign ICACHE_wdata[1] = 1'b0;
  assign ICACHE_wdata[2] = 1'b0;
  assign ICACHE_wdata[3] = 1'b0;
  assign ICACHE_wdata[4] = 1'b0;
  assign ICACHE_wdata[5] = 1'b0;
  assign ICACHE_wdata[6] = 1'b0;
  assign ICACHE_wdata[7] = 1'b0;
  assign ICACHE_wdata[8] = 1'b0;
  assign ICACHE_wdata[9] = 1'b0;
  assign ICACHE_wdata[10] = 1'b0;
  assign ICACHE_wdata[11] = 1'b0;
  assign ICACHE_wdata[12] = 1'b0;
  assign ICACHE_wdata[13] = 1'b0;
  assign ICACHE_wdata[14] = 1'b0;
  assign ICACHE_wdata[15] = 1'b0;
  assign ICACHE_wdata[16] = 1'b0;
  assign ICACHE_wdata[17] = 1'b0;
  assign ICACHE_wdata[18] = 1'b0;
  assign ICACHE_wdata[19] = 1'b0;
  assign ICACHE_wdata[20] = 1'b0;
  assign ICACHE_wdata[21] = 1'b0;
  assign ICACHE_wdata[22] = 1'b0;
  assign ICACHE_wdata[23] = 1'b0;
  assign ICACHE_wdata[24] = 1'b0;
  assign ICACHE_wdata[25] = 1'b0;
  assign ICACHE_wdata[26] = 1'b0;
  assign ICACHE_wdata[27] = 1'b0;
  assign ICACHE_wdata[28] = 1'b0;
  assign ICACHE_wdata[29] = 1'b0;
  assign ICACHE_wdata[30] = 1'b0;
  assign ICACHE_wdata[31] = 1'b0;
  assign ICACHE_wen = 1'b0;
  assign ICACHE_ren = 1'b1;

  BUFX4 U269 ( .A(Instruction[17]), .Y(n286) );
  BUFX4 U270 ( .A(Instruction[22]), .Y(n291) );
  OAI31X2 U271 ( .A0(n297), .A1(EX_MEM_RegisterRd[4]), .A2(
        EX_MEM_RegisterRd[3]), .B0(EX_MEM_WBControl[1]), .Y(n298) );
  CLKINVX8 U272 ( .A(EX_MEM_RegisterRd[3]), .Y(n314) );
  CLKINVX1 U273 ( .A(MEM_WB_RegisterRd[4]), .Y(n323) );
  OA21X2 U274 ( .A0(n242), .A1(MEM_WB_RegisterRd[3]), .B0(MEM_WB_WBControl[1]), 
        .Y(n327) );
  XOR2X1 U275 ( .A(n323), .B(ID_EX_RegisterRt[4]), .Y(n305) );
  XOR2X1 U276 ( .A(n315), .B(ID_EX_RegisterRt[4]), .Y(n304) );
  XOR2X1 U277 ( .A(n313), .B(ID_EX_RegisterRt[0]), .Y(n303) );
  CLKINVX1 U278 ( .A(EX_MEM_RegisterRd[2]), .Y(n311) );
  XOR2X1 U279 ( .A(n314), .B(ID_EX_RegisterRt[3]), .Y(n300) );
  INVX3 U280 ( .A(EX_MEM_RegisterRd[0]), .Y(n313) );
  XOR2X1 U281 ( .A(ID_EX_RegisterRt[1]), .B(n291), .Y(n81) );
  NOR2X4 U282 ( .A(n309), .B(n238), .Y(ForwardB[0]) );
  OR2X4 U283 ( .A(PredictMiss), .B(n276), .Y(IF_Flush) );
  CLKMX2X2 U284 ( .A(Buf_ALUresult[9]), .B(MemoryData[9]), .S0(n278), .Y(n269)
         );
  CLKINVX1 U285 ( .A(n74), .Y(n335) );
  CLKINVX1 U286 ( .A(EX_MEM_RegisterRd[4]), .Y(n315) );
  OR3XL U287 ( .A(n292), .B(n293), .C(n291), .Y(n204) );
  BUFX8 U288 ( .A(Instruction[19]), .Y(n288) );
  CLKBUFX3 U289 ( .A(Instruction[16]), .Y(n285) );
  CLKBUFX3 U290 ( .A(Instruction[21]), .Y(n290) );
  CLKBUFX6 U291 ( .A(Instruction[23]), .Y(n292) );
  BUFX4 U292 ( .A(Instruction[18]), .Y(n287) );
  BUFX4 U293 ( .A(Instruction[24]), .Y(n293) );
  CLKBUFX6 U294 ( .A(Instruction[25]), .Y(n294) );
  CLKBUFX6 U295 ( .A(Instruction[20]), .Y(n289) );
  BUFX2 U296 ( .A(needStall), .Y(n295) );
  XNOR2X1 U297 ( .A(MEM_WB_RegisterRd[1]), .B(ID_EX_RegisterRt[1]), .Y(n237)
         );
  OR3X2 U298 ( .A(n306), .B(n308), .C(n307), .Y(n238) );
  CLKINVX1 U299 ( .A(EX_MEM_RegisterRd[1]), .Y(n312) );
  NAND3BX1 U300 ( .AN(EX_MEM_RegisterRd[1]), .B(n313), .C(n311), .Y(n297) );
  BUFX12 U301 ( .A(N199), .Y(DCACHE_ren) );
  NOR2BX1 U302 ( .AN(EX_MEM_MEMControl[1]), .B(EX_MEM_MEMControl[0]), .Y(N199)
         );
  BUFX12 U303 ( .A(N202), .Y(DCACHE_wen) );
  NOR2BX1 U304 ( .AN(EX_MEM_MEMControl[0]), .B(EX_MEM_MEMControl[1]), .Y(N202)
         );
  OR4X1 U305 ( .A(MEM_WB_RegisterRd[4]), .B(MEM_WB_RegisterRd[1]), .C(
        MEM_WB_RegisterRd[0]), .D(MEM_WB_RegisterRd[2]), .Y(n242) );
  MX2X1 U306 ( .A(Buf_ALUresult[4]), .B(MemoryData[4]), .S0(n278), .Y(n266) );
  INVX4 U307 ( .A(n298), .Y(n322) );
  AND3X4 U308 ( .A(n301), .B(n300), .C(n299), .Y(n302) );
  MX2XL U309 ( .A(Buf_ALUresult[13]), .B(MemoryData[13]), .S0(n279), .Y(n272)
         );
  INVXL U310 ( .A(MEM_WB_RegisterRd[1]), .Y(n324) );
  NAND4X6 U311 ( .A(n322), .B(n304), .C(n303), .D(n302), .Y(n310) );
  CLKMX2X2 U312 ( .A(PCbranched[25]), .B(next_ReadData1[25]), .S0(n276), .Y(
        PCJump_JRChecked[25]) );
  NAND4X4 U313 ( .A(n327), .B(n310), .C(n305), .D(n237), .Y(n309) );
  XOR2XL U314 ( .A(n312), .B(ID_EX_RegisterRt[1]), .Y(n301) );
  AO22X1 U315 ( .A0(PCbranched[15]), .A1(n75), .B0(next_ReadData1[15]), .B1(
        n277), .Y(PCJump_JRChecked[15]) );
  XOR2XL U316 ( .A(n311), .B(ID_EX_RegisterRt[2]), .Y(n299) );
  MX2XL U317 ( .A(Buf_ALUresult[20]), .B(MemoryData[20]), .S0(n279), .Y(n250)
         );
  MX2X1 U318 ( .A(Buf_ALUresult[24]), .B(MemoryData[24]), .S0(n279), .Y(n254)
         );
  AO22X1 U319 ( .A0(PCbranched[21]), .A1(n75), .B0(next_ReadData1[21]), .B1(
        n277), .Y(PCJump_JRChecked[21]) );
  AO22X1 U320 ( .A0(PCbranched[9]), .A1(n75), .B0(next_ReadData1[9]), .B1(n276), .Y(PCJump_JRChecked[9]) );
  AO22X1 U321 ( .A0(PCbranched[5]), .A1(n75), .B0(next_ReadData1[5]), .B1(n277), .Y(PCJump_JRChecked[5]) );
  MX2XL U322 ( .A(Buf_ALUresult[0]), .B(MemoryData[0]), .S0(n278), .Y(n262) );
  MX2XL U323 ( .A(Buf_ALUresult[11]), .B(MemoryData[11]), .S0(n278), .Y(n243)
         );
  AO22X2 U324 ( .A0(PCbranched[17]), .A1(n275), .B0(next_ReadData1[17]), .B1(
        n277), .Y(PCJump_JRChecked[17]) );
  AO22X2 U325 ( .A0(PCbranched[23]), .A1(n275), .B0(next_ReadData1[23]), .B1(
        n277), .Y(PCJump_JRChecked[23]) );
  OA21XL U326 ( .A0(n127), .A1(n128), .B0(Branch), .Y(BrForwardB[1]) );
  OA21XL U327 ( .A0(n155), .A1(n156), .B0(Branch), .Y(BrForwardA[1]) );
  OA21XL U328 ( .A0(n129), .A1(n128), .B0(Branch), .Y(BrForwardB[0]) );
  OA21XL U329 ( .A0(n157), .A1(n156), .B0(Branch), .Y(BrForwardA[0]) );
  CLKINVX1 U330 ( .A(n73), .Y(n333) );
  NAND4XL U331 ( .A(n322), .B(n321), .C(n320), .D(n319), .Y(n332) );
  XOR2XL U332 ( .A(n312), .B(ID_EX_RegisterRs[1]), .Y(n320) );
  XOR2XL U333 ( .A(n311), .B(ID_EX_RegisterRs[2]), .Y(n321) );
  XOR2XL U334 ( .A(n315), .B(ID_EX_RegisterRs[4]), .Y(n316) );
  XOR2XL U335 ( .A(n313), .B(ID_EX_RegisterRs[0]), .Y(n318) );
  XOR2XL U336 ( .A(n314), .B(ID_EX_RegisterRs[3]), .Y(n317) );
  MX2X1 U337 ( .A(Buf_ALUresult[14]), .B(MemoryData[14]), .S0(n279), .Y(n274)
         );
  MX2X1 U338 ( .A(Buf_ALUresult[1]), .B(MemoryData[1]), .S0(n278), .Y(n261) );
  MX2XL U339 ( .A(Buf_ALUresult[16]), .B(MemoryData[16]), .S0(n279), .Y(n246)
         );
  XOR2XL U340 ( .A(n287), .B(ID_EX_RegisterRd[2]), .Y(n151) );
  XOR2XL U341 ( .A(n292), .B(ID_EX_RegisterRd[2]), .Y(n180) );
  XOR2XL U342 ( .A(n288), .B(ID_EX_RegisterRd[3]), .Y(n152) );
  XOR2XL U343 ( .A(n293), .B(ID_EX_RegisterRd[3]), .Y(n181) );
  XNOR2XL U344 ( .A(ID_EX_RegisterRd[1]), .B(n286), .Y(n148) );
  XNOR2XL U345 ( .A(ID_EX_RegisterRd[1]), .B(n291), .Y(n177) );
  NOR3XL U346 ( .A(n91), .B(Instruction[28]), .C(n353), .Y(Jump) );
  MX2XL U347 ( .A(Buf_ALUresult[18]), .B(MemoryData[18]), .S0(n279), .Y(n248)
         );
  MX2XL U348 ( .A(Buf_ALUresult[22]), .B(MemoryData[22]), .S0(n279), .Y(n252)
         );
  MX2XL U349 ( .A(Buf_ALUresult[23]), .B(MemoryData[23]), .S0(n279), .Y(n251)
         );
  MX2XL U350 ( .A(Buf_ALUresult[19]), .B(MemoryData[19]), .S0(n279), .Y(n247)
         );
  MX2XL U351 ( .A(Buf_ALUresult[21]), .B(MemoryData[21]), .S0(n279), .Y(n249)
         );
  MX2XL U352 ( .A(Buf_ALUresult[17]), .B(MemoryData[17]), .S0(n279), .Y(n245)
         );
  MX2X1 U353 ( .A(Buf_ALUresult[26]), .B(MemoryData[26]), .S0(n279), .Y(n256)
         );
  MX2XL U354 ( .A(Buf_ALUresult[27]), .B(MemoryData[27]), .S0(n279), .Y(n255)
         );
  MX2XL U355 ( .A(Buf_ALUresult[31]), .B(MemoryData[31]), .S0(n279), .Y(n259)
         );
  MX2XL U356 ( .A(Buf_ALUresult[30]), .B(MemoryData[30]), .S0(n279), .Y(n260)
         );
  MX2XL U357 ( .A(Buf_ALUresult[29]), .B(MemoryData[29]), .S0(n279), .Y(n257)
         );
  MX2XL U358 ( .A(Buf_ALUresult[28]), .B(MemoryData[28]), .S0(n278), .Y(n258)
         );
  AOI211XL U359 ( .A0(n77), .A1(n345), .B0(n153), .C0(n344), .Y(n144) );
  AOI211XL U360 ( .A0(n80), .A1(n345), .B0(n182), .C0(n344), .Y(n173) );
  XOR2XL U361 ( .A(MEM_WB_RegisterRd[3]), .B(n288), .Y(n140) );
  XOR2XL U362 ( .A(MEM_WB_RegisterRd[3]), .B(n293), .Y(n169) );
  NOR3XL U363 ( .A(Instruction[26]), .B(Instruction[27]), .C(n91), .Y(n159) );
  INVX1 U364 ( .A(Instruction[28]), .Y(n352) );
  INVX1 U365 ( .A(Instruction[27]), .Y(n353) );
  INVX1 U366 ( .A(Instruction[29]), .Y(n350) );
  INVXL U367 ( .A(Instruction[30]), .Y(n349) );
  XNOR2XL U368 ( .A(EX_MEM_RegisterRd[1]), .B(n286), .Y(n134) );
  XNOR2XL U369 ( .A(EX_MEM_RegisterRd[0]), .B(n285), .Y(n136) );
  XNOR2XL U370 ( .A(EX_MEM_RegisterRd[4]), .B(n289), .Y(n135) );
  XNOR2XL U371 ( .A(EX_MEM_RegisterRd[1]), .B(n291), .Y(n163) );
  XNOR2XL U372 ( .A(EX_MEM_RegisterRd[4]), .B(n294), .Y(n164) );
  XNOR2XL U373 ( .A(EX_MEM_RegisterRd[0]), .B(n290), .Y(n165) );
  XOR2XL U374 ( .A(MEM_WB_RegisterRd[4]), .B(n289), .Y(n143) );
  XOR2XL U375 ( .A(MEM_WB_RegisterRd[4]), .B(n294), .Y(n172) );
  XOR2XL U376 ( .A(n287), .B(EX_MEM_RegisterRd[2]), .Y(n138) );
  XOR2XL U377 ( .A(n288), .B(EX_MEM_RegisterRd[3]), .Y(n139) );
  XOR2XL U378 ( .A(n292), .B(EX_MEM_RegisterRd[2]), .Y(n167) );
  XOR2XL U379 ( .A(n293), .B(EX_MEM_RegisterRd[3]), .Y(n168) );
  XOR2XL U380 ( .A(n285), .B(ID_EX_RegisterRd[0]), .Y(n146) );
  XOR2XL U381 ( .A(n290), .B(ID_EX_RegisterRd[0]), .Y(n175) );
  XOR2XL U382 ( .A(MEM_WB_RegisterRd[0]), .B(n290), .Y(n171) );
  XOR2XL U383 ( .A(MEM_WB_RegisterRd[0]), .B(n285), .Y(n142) );
  XOR2XL U384 ( .A(MEM_WB_RegisterRd[1]), .B(n286), .Y(n141) );
  XOR2XL U385 ( .A(MEM_WB_RegisterRd[1]), .B(n291), .Y(n170) );
  XOR2XL U386 ( .A(MEM_WB_RegisterRd[2]), .B(n292), .Y(n162) );
  XOR2XL U387 ( .A(MEM_WB_RegisterRd[2]), .B(n287), .Y(n133) );
  INVXL U388 ( .A(Instruction[31]), .Y(n347) );
  XNOR2XL U389 ( .A(ID_EX_RegisterRd[4]), .B(n289), .Y(n154) );
  XNOR2XL U390 ( .A(ID_EX_RegisterRd[4]), .B(n294), .Y(n183) );
  INVXL U391 ( .A(EX_MEM_WBControl[1]), .Y(n343) );
  INVXL U392 ( .A(MEM_WB_WBControl[1]), .Y(n342) );
  NOR3XL U393 ( .A(n294), .B(Instruction[6]), .C(Instruction[3]), .Y(n196) );
  NOR4XL U394 ( .A(n204), .B(n288), .C(n290), .D(n289), .Y(n198) );
  NOR3XL U395 ( .A(Instruction[30]), .B(Instruction[31]), .C(n350), .Y(n192)
         );
  OAI31XL U396 ( .A0(n348), .A1(n352), .A2(n353), .B0(n191), .Y(n189) );
  NAND4XL U397 ( .A(n192), .B(Instruction[26]), .C(Instruction[28]), .D(n353), 
        .Y(n191) );
  AOI2BB2XL U398 ( .B0(Instruction[27]), .B1(n347), .A0N(n348), .A1N(n352), 
        .Y(n193) );
  NAND2XL U399 ( .A(n188), .B(Instruction[27]), .Y(n184) );
  NAND2XL U400 ( .A(Instruction[26]), .B(n352), .Y(n195) );
  NAND4XL U401 ( .A(Instruction[31]), .B(Instruction[27]), .C(n186), .D(n351), 
        .Y(n89) );
  NOR2XL U402 ( .A(Instruction[30]), .B(Instruction[29]), .Y(n186) );
  NAND4XL U403 ( .A(n351), .B(n349), .C(Instruction[27]), .D(n187), .Y(n90) );
  XOR2XL U404 ( .A(ID_EX_RegisterRt[2]), .B(MEM_WB_RegisterRd[2]), .Y(n308) );
  XOR2XL U405 ( .A(ID_EX_RegisterRt[0]), .B(MEM_WB_RegisterRd[0]), .Y(n307) );
  XOR2XL U406 ( .A(ID_EX_RegisterRt[3]), .B(MEM_WB_RegisterRd[3]), .Y(n306) );
  INVX3 U407 ( .A(n275), .Y(n276) );
  INVX3 U408 ( .A(n275), .Y(n277) );
  CLKINVX1 U409 ( .A(n185), .Y(n55) );
  CLKINVX1 U410 ( .A(n310), .Y(ForwardB[1]) );
  AO22X1 U411 ( .A0(PCbranched[6]), .A1(n275), .B0(next_ReadData1[6]), .B1(
        n277), .Y(PCJump_JRChecked[6]) );
  CLKMX2X2 U412 ( .A(PCbranched[27]), .B(next_ReadData1[27]), .S0(n276), .Y(
        PCJump_JRChecked[27]) );
  AO22X1 U413 ( .A0(PCbranched[11]), .A1(n275), .B0(next_ReadData1[11]), .B1(
        n276), .Y(PCJump_JRChecked[11]) );
  CLKMX2X2 U414 ( .A(PCbranched[29]), .B(next_ReadData1[29]), .S0(n276), .Y(
        PCJump_JRChecked[29]) );
  CLKMX2X2 U415 ( .A(PCbranched[28]), .B(next_ReadData1[28]), .S0(n276), .Y(
        PCJump_JRChecked[28]) );
  AO22X1 U416 ( .A0(PCbranched[16]), .A1(n275), .B0(next_ReadData1[16]), .B1(
        n277), .Y(PCJump_JRChecked[16]) );
  AO22X1 U417 ( .A0(PCbranched[18]), .A1(n275), .B0(next_ReadData1[18]), .B1(
        n277), .Y(PCJump_JRChecked[18]) );
  AO22X1 U418 ( .A0(PCbranched[19]), .A1(n275), .B0(next_ReadData1[19]), .B1(
        n277), .Y(PCJump_JRChecked[19]) );
  AO22X1 U419 ( .A0(PCbranched[20]), .A1(n275), .B0(next_ReadData1[20]), .B1(
        n277), .Y(PCJump_JRChecked[20]) );
  AO22X1 U420 ( .A0(PCbranched[22]), .A1(n275), .B0(next_ReadData1[22]), .B1(
        n277), .Y(PCJump_JRChecked[22]) );
  AO22X1 U421 ( .A0(PCbranched[24]), .A1(n275), .B0(next_ReadData1[24]), .B1(
        n277), .Y(PCJump_JRChecked[24]) );
  AO22X1 U422 ( .A0(PCbranched[8]), .A1(n75), .B0(next_ReadData1[8]), .B1(n277), .Y(PCJump_JRChecked[8]) );
  AO22X1 U423 ( .A0(PCbranched[10]), .A1(n275), .B0(next_ReadData1[10]), .B1(
        n276), .Y(PCJump_JRChecked[10]) );
  AO22X1 U424 ( .A0(PCbranched[12]), .A1(n275), .B0(next_ReadData1[12]), .B1(
        n276), .Y(PCJump_JRChecked[12]) );
  AO22X1 U425 ( .A0(PCbranched[14]), .A1(n275), .B0(next_ReadData1[14]), .B1(
        n276), .Y(PCJump_JRChecked[14]) );
  AO22X1 U426 ( .A0(PCbranched[7]), .A1(n275), .B0(next_ReadData1[7]), .B1(
        n277), .Y(PCJump_JRChecked[7]) );
  AO22X1 U427 ( .A0(PCbranched[13]), .A1(n275), .B0(next_ReadData1[13]), .B1(
        n276), .Y(PCJump_JRChecked[13]) );
  CLKMX2X2 U428 ( .A(PCbranched[26]), .B(next_ReadData1[26]), .S0(n276), .Y(
        PCJump_JRChecked[26]) );
  CLKINVX1 U429 ( .A(n332), .Y(ForwardA[1]) );
  NAND3X1 U430 ( .A(n349), .B(n347), .C(n350), .Y(n91) );
  CLKBUFX3 U431 ( .A(MEM_WB_WBControl[0]), .Y(n278) );
  CLKBUFX3 U432 ( .A(MEM_WB_WBControl[0]), .Y(n279) );
  AO22X1 U433 ( .A0(PCbranched[2]), .A1(n275), .B0(next_ReadData1[2]), .B1(
        n277), .Y(PCJump_JRChecked[2]) );
  AO22X1 U434 ( .A0(PCbranched[3]), .A1(n275), .B0(next_ReadData1[3]), .B1(
        n277), .Y(PCJump_JRChecked[3]) );
  NOR2BX2 U435 ( .AN(n159), .B(n352), .Y(Branch) );
  NOR2X1 U436 ( .A(n129), .B(n130), .Y(n127) );
  NOR2X1 U437 ( .A(n157), .B(n158), .Y(n155) );
  AOI21X1 U438 ( .A0(n353), .A1(n188), .B0(n189), .Y(n185) );
  AOI21X1 U439 ( .A0(n335), .A1(n334), .B0(n333), .Y(n241) );
  NAND2X1 U440 ( .A(n159), .B(n352), .Y(n190) );
  CLKINVX1 U441 ( .A(n189), .Y(n334) );
  NAND2X1 U442 ( .A(n190), .B(n184), .Y(n74) );
  CLKINVX1 U443 ( .A(n188), .Y(n348) );
  CLKBUFX3 U444 ( .A(n75), .Y(n275) );
  CLKINVX1 U445 ( .A(n195), .Y(n351) );
  OR3X2 U446 ( .A(n286), .B(n287), .C(n285), .Y(n202) );
  CLKINVX1 U447 ( .A(n89), .Y(n57) );
  AO22X1 U448 ( .A0(PCbranched[4]), .A1(n75), .B0(next_ReadData1[4]), .B1(n277), .Y(PCJump_JRChecked[4]) );
  AO22X1 U449 ( .A0(PCbranched[0]), .A1(n275), .B0(next_ReadData1[0]), .B1(
        n276), .Y(PCJump_JRChecked[0]) );
  AO22X1 U450 ( .A0(PCbranched[1]), .A1(n275), .B0(next_ReadData1[1]), .B1(
        n277), .Y(PCJump_JRChecked[1]) );
  CLKMX2X2 U451 ( .A(PCbranched[31]), .B(next_ReadData1[31]), .S0(n276), .Y(
        PCJump_JRChecked[31]) );
  CLKMX2X2 U452 ( .A(PCbranched[30]), .B(next_ReadData1[30]), .S0(n276), .Y(
        PCJump_JRChecked[30]) );
  NOR4X1 U453 ( .A(n331), .B(n330), .C(n329), .D(n328), .Y(ForwardA[0]) );
  XOR2X1 U454 ( .A(ID_EX_RegisterRs[2]), .B(MEM_WB_RegisterRd[2]), .Y(n330) );
  XOR2X1 U455 ( .A(ID_EX_RegisterRs[3]), .B(MEM_WB_RegisterRd[3]), .Y(n328) );
  XOR2X1 U456 ( .A(ID_EX_RegisterRs[0]), .B(MEM_WB_RegisterRd[0]), .Y(n329) );
  AND3X2 U457 ( .A(n318), .B(n317), .C(n316), .Y(n319) );
  NAND4X1 U458 ( .A(n327), .B(n332), .C(n326), .D(n325), .Y(n331) );
  XOR2X1 U459 ( .A(n323), .B(ID_EX_RegisterRs[4]), .Y(n326) );
  XOR2X1 U460 ( .A(n324), .B(ID_EX_RegisterRs[1]), .Y(n325) );
  CLKMX2X2 U461 ( .A(Buf_ALUresult[15]), .B(MemoryData[15]), .S0(n279), .Y(
        n244) );
  XOR2X1 U462 ( .A(ID_EX_RegisterRt[3]), .B(Instruction[19]), .Y(n87) );
  XOR2X1 U463 ( .A(ID_EX_RegisterRt[3]), .B(Instruction[24]), .Y(n84) );
  XOR2X1 U464 ( .A(ID_EX_RegisterRt[2]), .B(Instruction[23]), .Y(n85) );
  XOR2X1 U465 ( .A(ID_EX_RegisterRt[2]), .B(Instruction[18]), .Y(n88) );
  XOR2X1 U466 ( .A(ID_EX_RegisterRt[4]), .B(Instruction[25]), .Y(n80) );
  XOR2X1 U467 ( .A(ID_EX_RegisterRt[4]), .B(Instruction[20]), .Y(n77) );
  XOR2X1 U468 ( .A(ID_EX_RegisterRt[1]), .B(n286), .Y(n78) );
  XOR2X1 U469 ( .A(ID_EX_RegisterRt[0]), .B(n290), .Y(n83) );
  XOR2X1 U470 ( .A(ID_EX_RegisterRt[0]), .B(n285), .Y(n86) );
  CLKMX2X2 U471 ( .A(Buf_ALUresult[25]), .B(MemoryData[25]), .S0(n279), .Y(
        n253) );
  CLKMX2X2 U472 ( .A(Buf_ALUresult[3]), .B(MemoryData[3]), .S0(n278), .Y(n263)
         );
  CLKMX2X2 U473 ( .A(Buf_ALUresult[2]), .B(MemoryData[2]), .S0(n278), .Y(n264)
         );
  CLKMX2X2 U474 ( .A(Buf_ALUresult[5]), .B(MemoryData[5]), .S0(n278), .Y(n265)
         );
  CLKMX2X2 U475 ( .A(Buf_ALUresult[7]), .B(MemoryData[7]), .S0(n278), .Y(n267)
         );
  CLKMX2X2 U476 ( .A(Buf_ALUresult[6]), .B(MemoryData[6]), .S0(n278), .Y(n268)
         );
  CLKMX2X2 U477 ( .A(Buf_ALUresult[8]), .B(MemoryData[8]), .S0(n278), .Y(n270)
         );
  CLKMX2X2 U478 ( .A(Buf_ALUresult[10]), .B(MemoryData[10]), .S0(n278), .Y(
        n271) );
  CLKMX2X2 U479 ( .A(Buf_ALUresult[12]), .B(MemoryData[12]), .S0(n279), .Y(
        n273) );
  AND2X2 U480 ( .A(ID_EX_MEMControl[1]), .B(n76), .Y(N182) );
  OAI33X1 U481 ( .A0(n77), .A1(n78), .A2(n79), .B0(n80), .B1(n81), .B2(n82), 
        .Y(n76) );
  OR3X2 U482 ( .A(n86), .B(n87), .C(n88), .Y(n79) );
  OR3X2 U483 ( .A(n83), .B(n84), .C(n85), .Y(n82) );
  OR2X1 U484 ( .A(DCACHE_stall), .B(ICACHE_stall), .Y(needStall) );
  CLKBUFX3 U485 ( .A(Immediate_SE[8]), .Y(n282) );
  CLKBUFX3 U486 ( .A(Immediate_SE[7]), .Y(n281) );
  CLKBUFX3 U487 ( .A(Immediate_SE[9]), .Y(n283) );
  CLKBUFX3 U488 ( .A(Immediate_SE[6]), .Y(n280) );
  CLKBUFX3 U489 ( .A(Immediate_SE[10]), .Y(n284) );
  OAI211X1 U490 ( .A0(n148), .A1(n345), .B0(n149), .C0(n150), .Y(n147) );
  OAI21XL U491 ( .A0(n151), .A1(n152), .B0(ID_EX_EXControl[4]), .Y(n149) );
  OAI21XL U492 ( .A0(n87), .A1(n88), .B0(n345), .Y(n150) );
  OAI211X1 U493 ( .A0(n177), .A1(n345), .B0(n178), .C0(n179), .Y(n176) );
  OAI21XL U494 ( .A0(n180), .A1(n181), .B0(ID_EX_EXControl[4]), .Y(n178) );
  OAI21XL U495 ( .A0(n84), .A1(n85), .B0(n345), .Y(n179) );
  NAND4X1 U496 ( .A(n134), .B(n135), .C(n136), .D(n137), .Y(n130) );
  NAND4X1 U497 ( .A(n163), .B(n164), .C(n165), .D(n166), .Y(n158) );
  INVX3 U498 ( .A(ID_EX_EXControl[4]), .Y(n345) );
  NOR3X1 U499 ( .A(n138), .B(n343), .C(n139), .Y(n137) );
  NOR3X1 U500 ( .A(n167), .B(n343), .C(n168), .Y(n166) );
  AND2X2 U501 ( .A(n144), .B(n145), .Y(n129) );
  AOI221XL U502 ( .A0(n78), .A1(n345), .B0(ID_EX_EXControl[4]), .B1(n146), 
        .C0(n147), .Y(n145) );
  OAI2BB2XL U503 ( .B0(n154), .B1(n345), .A0N(n345), .A1N(n86), .Y(n153) );
  AND2X2 U504 ( .A(n173), .B(n174), .Y(n157) );
  AOI221XL U505 ( .A0(n81), .A1(n345), .B0(ID_EX_EXControl[4]), .B1(n175), 
        .C0(n176), .Y(n174) );
  OAI2BB2XL U506 ( .B0(n183), .B1(n345), .A0N(n345), .A1N(n83), .Y(n182) );
  CLKINVX1 U507 ( .A(ID_EX_WBControl[1]), .Y(n344) );
  AND2X2 U508 ( .A(n131), .B(n132), .Y(n128) );
  NOR4X1 U509 ( .A(n140), .B(n141), .C(n142), .D(n143), .Y(n131) );
  NOR4BX1 U510 ( .AN(n130), .B(n129), .C(n342), .D(n133), .Y(n132) );
  AND2X2 U511 ( .A(n160), .B(n161), .Y(n156) );
  NOR4X1 U512 ( .A(n169), .B(n170), .C(n171), .D(n172), .Y(n160) );
  NOR4BX1 U513 ( .AN(n158), .B(n157), .C(n342), .D(n162), .Y(n161) );
  NAND3BX1 U514 ( .AN(\ALUOp[0] ), .B(n241), .C(n340), .Y(n75) );
  AND3X2 U515 ( .A(Instruction[3]), .B(n185), .C(n341), .Y(n340) );
  NOR2BX1 U516 ( .AN(n192), .B(Instruction[26]), .Y(n188) );
  NAND4X1 U517 ( .A(n196), .B(n197), .C(n198), .D(n199), .Y(n73) );
  NOR3X1 U518 ( .A(Instruction[7]), .B(Instruction[9]), .C(Instruction[8]), 
        .Y(n197) );
  NAND4X1 U519 ( .A(n73), .B(n349), .C(n193), .D(n194), .Y(\ALUOp[0] ) );
  AOI222XL U520 ( .A0(Instruction[31]), .A1(n195), .B0(Instruction[28]), .B1(
        n350), .C0(n351), .C1(n353), .Y(n194) );
  AND4X1 U521 ( .A(n341), .B(n346), .C(n200), .D(n201), .Y(n199) );
  NOR3X1 U522 ( .A(Instruction[10]), .B(Instruction[12]), .C(Instruction[11]), 
        .Y(n200) );
  NOR4X1 U523 ( .A(n202), .B(Instruction[13]), .C(Instruction[15]), .D(
        Instruction[14]), .Y(n201) );
  CLKINVX1 U524 ( .A(n190), .Y(n346) );
  CLKINVX1 U525 ( .A(n339), .Y(n341) );
  NAND4BX1 U526 ( .AN(n203), .B(n338), .C(n337), .D(n336), .Y(n339) );
  CLKINVX1 U527 ( .A(Instruction[0]), .Y(n337) );
  CLKINVX1 U528 ( .A(Instruction[1]), .Y(n336) );
  CLKINVX1 U529 ( .A(Instruction[2]), .Y(n338) );
  NAND4X1 U530 ( .A(n184), .B(n185), .C(n90), .D(n89), .Y(ALUSrc) );
  CLKINVX1 U531 ( .A(n90), .Y(n56) );
  CLKINVX1 U532 ( .A(n72), .Y(n54) );
  AOI211X1 U533 ( .A0(n73), .A1(n74), .B0(n55), .C0(n57), .Y(n72) );
  OR2X1 U534 ( .A(Instruction[5]), .B(Instruction[4]), .Y(n203) );
  NOR2X1 U535 ( .A(n347), .B(n350), .Y(n187) );
  CLKBUFX3 U536 ( .A(rst), .Y(n296) );
  InstructionFetch_test_1 IF ( .clk(clk), .rst(n296), .stall(n295), .PCWrite(
        N182), .PCJumpJRorBranch(PCJump_JRChecked), .IF_ID_Write(N182), 
        .IF_Flush(IF_Flush), .PCadd4(PCadd4), .Instruction(Instruction), .PC(
        ICACHE_addr), .read_Instruction(ICACHE_rdata), .PredictMiss(
        PredictMiss), .BranchTaken(BranchTaken), .PCBuffer_valid(
        PCBuffer_valid), .test_si(n3), .test_so(test_so), .test_se(test_se) );
  InstructionDecode_test_1 ID ( .clk(clk), .rst(n296), .stall(n295), .PCadd4(
        PCadd4), .Instruction({Instruction[31:26], n294, n293, n292, n291, 
        n290, n289, n288, n287, n286, n285, Instruction[15:0]}), .PCbranched(
        PCbranched), .Reg_W(MEM_WB_RegisterRd), .WriteData({n259, n260, n257, 
        n258, n255, n256, n253, n254, n251, n252, n249, n250, n247, n248, n245, 
        n246, n244, n274, n272, n273, n243, n271, n269, n270, n267, n268, n265, 
        n266, n263, n264, n261, n262}), .WB(ID_EX_WBControl), .MEM({
        SYNOPSYS_UNCONNECTED__0, ID_EX_MEMControl[1:0]}), .EX(ID_EX_EXControl), 
        .RData1(ReadData1), .RData2(ReadData2), .next_RData1(next_ReadData1), 
        .Immediate_SE(Immediate_SE), .RegisterRd(ID_EX_RegisterRd), 
        .RegisterRs(ID_EX_RegisterRs), .RegisterRt(ID_EX_RegisterRt), 
        .MEM_RegWrite(MEM_WB_WBControl[1]), .RegDst(n346), .Jump(Jump), 
        .Branch(Branch), .MemRead(n57), .MemtoReg(n57), .MemWrite(n56), 
        .ALUOp({n55, n241, \ALUOp[0] }), .ALUSrc(ALUSrc), .RegWrite(n54), 
        .Bubble(N182), .PCBuffer_valid(PCBuffer_valid), .EX_RegWriteData(
        next_ALUresult), .MEM_RegWriteData(DCACHE_addr), .BrForwardA(
        BrForwardA), .BrForwardB(BrForwardB), .PredictMiss(PredictMiss), 
        .BranchTaken(BranchTaken), .test_si2(n4), .test_si1(test_si), 
        .test_so2(n3), .test_so1(n6), .test_se(test_se) );
  Execution_test_1 EX ( .clk(clk), .rst(n296), .stall(n295), .ID_WB(
        ID_EX_WBControl), .ID_MEM({1'b0, ID_EX_MEMControl[1:0]}), .ID_EX(
        ID_EX_EXControl), .RData1(ReadData1), .RData2(ReadData2), 
        .Immediate_SE({Immediate_SE[31:11], n284, n283, n282, n281, n280, 
        Immediate_SE[5:0]}), .ID_RegisterRt(ID_EX_RegisterRt), .ID_RegisterRd(
        ID_EX_RegisterRd), .WB(EX_MEM_WBControl), .MEM(EX_MEM_MEMControl), 
        .next_ALUresult(next_ALUresult), .ALUresult(DCACHE_addr), 
        .MEMWriteData(DCACHE_wdata), .RegisterRd(EX_MEM_RegisterRd), .WBData({
        n259, n260, n257, n258, n255, n256, n253, n254, n251, n252, n249, n250, 
        n247, n248, n245, n246, n244, n274, n272, n273, n243, n271, n269, n270, 
        n267, n268, n265, n266, n263, n264, n261, n262}), .ForwardA(ForwardA), 
        .ForwardB(ForwardB), .test_si(n5), .test_so(n4), .test_se(test_se) );
  DataMemory_test_1 DMEM ( .clk(clk), .rst(n296), .stall(n295), .EX_WB(
        EX_MEM_WBControl), .EX_MEM(EX_MEM_MEMControl), .EX_ALUresult(
        DCACHE_addr), .EX_RegisterRd(EX_MEM_RegisterRd), .MEMWriteData(
        DCACHE_wdata), .WB(MEM_WB_WBControl), .MemoryData(MemoryData), 
        .ALUresult(Buf_ALUresult), .RegisterRd(MEM_WB_RegisterRd), 
        .read_MemoryData(DCACHE_rdata), .test_si(n6), .test_so(n5), .test_se(
        test_se) );
endmodule

module CHIP ( 	clk, rst, ICACHE_addr, ICACHE_rdata, ICACHE_ren, 
				ICACHE_wen, ICACHE_wdata, ICACHE_stall, DCACHE_addr, DCACHE_rdata, 
				DCACHE_ren, DCACHE_wen, DCACHE_wdata, DCACHE_stall, test_si, test_so, 
				test_se );
				
		output [31:0] ICACHE_addr;
		input [31:0] ICACHE_rdata;
		output [31:0] ICACHE_wdata;
		output [31:0] DCACHE_addr;
		input [31:0] DCACHE_rdata;
		output [31:0] DCACHE_wdata;
		input clk, rst, ICACHE_stall, DCACHE_stall, test_si, test_se;
		output ICACHE_ren, ICACHE_wen, DCACHE_ren, DCACHE_wen, test_so;
		
		wire [31:0] ICACHE_addr_i;
		wire [31:0] ICACHE_rdata_i;
		wire [31:0] ICACHE_wdata_i;
		wire [31:0] DCACHE_addr_i;
		wire [31:0] DCACHE_rdata_i;
		wire [31:0] DCACHE_wdata_i;
		wire clk_i, rst_i, ICACHE_stall_i, DCACHE_stall_i, test_si_i, test_se_i;
		wire ICACHE_ren_i, ICACHE_wen_i, DCACHE_ren_i, DCACHE_wen_i, test_so_i;
		
		PDIDGZ ipad_clk (.PAD(clk), .C(clk_i));
		PDIDGZ ipad_rst (.PAD(rst), .C(rst_i));
		PDIDGZ ipad_ICACHE_stall (.PAD(ICACHE_stall), .C(ICACHE_stall_i));
		PDIDGZ ipad_DCACHE_stall (.PAD(DCACHE_stall), .C(DCACHE_stall_i));
		PDIDGZ ipad_test_si (.PAD(test_si), .C(test_si_i));
		PDIDGZ ipad_test_se (.PAD(test_se), .C(test_se_i));
		
		PDIDGZ ipad_ICACHE_rdata0 (.PAD(ICACHE_rdata[0]), .C(ICACHE_rdata_i[0]));
		PDIDGZ ipad_ICACHE_rdata1 (.PAD(ICACHE_rdata[1]), .C(ICACHE_rdata_i[1]));
		PDIDGZ ipad_ICACHE_rdata2 (.PAD(ICACHE_rdata[2]), .C(ICACHE_rdata_i[2]));
		PDIDGZ ipad_ICACHE_rdata3 (.PAD(ICACHE_rdata[3]), .C(ICACHE_rdata_i[3]));
		PDIDGZ ipad_ICACHE_rdata4 (.PAD(ICACHE_rdata[4]), .C(ICACHE_rdata_i[4]));
		PDIDGZ ipad_ICACHE_rdata5 (.PAD(ICACHE_rdata[5]), .C(ICACHE_rdata_i[5]));
		PDIDGZ ipad_ICACHE_rdata6 (.PAD(ICACHE_rdata[6]), .C(ICACHE_rdata_i[6]));
		PDIDGZ ipad_ICACHE_rdata7 (.PAD(ICACHE_rdata[7]), .C(ICACHE_rdata_i[7]));
		PDIDGZ ipad_ICACHE_rdata8 (.PAD(ICACHE_rdata[8]), .C(ICACHE_rdata_i[8]));
		PDIDGZ ipad_ICACHE_rdata9 (.PAD(ICACHE_rdata[9]), .C(ICACHE_rdata_i[9]));
		PDIDGZ ipad_ICACHE_rdata10 (.PAD(ICACHE_rdata[10]), .C(ICACHE_rdata_i[10]));
		PDIDGZ ipad_ICACHE_rdata11 (.PAD(ICACHE_rdata[11]), .C(ICACHE_rdata_i[11]));
		PDIDGZ ipad_ICACHE_rdata12 (.PAD(ICACHE_rdata[12]), .C(ICACHE_rdata_i[12]));
		PDIDGZ ipad_ICACHE_rdata13 (.PAD(ICACHE_rdata[13]), .C(ICACHE_rdata_i[13]));
		PDIDGZ ipad_ICACHE_rdata14 (.PAD(ICACHE_rdata[14]), .C(ICACHE_rdata_i[14]));
		PDIDGZ ipad_ICACHE_rdata15 (.PAD(ICACHE_rdata[15]), .C(ICACHE_rdata_i[15]));
		PDIDGZ ipad_ICACHE_rdata16 (.PAD(ICACHE_rdata[16]), .C(ICACHE_rdata_i[16]));
		PDIDGZ ipad_ICACHE_rdata17 (.PAD(ICACHE_rdata[17]), .C(ICACHE_rdata_i[17]));
		PDIDGZ ipad_ICACHE_rdata18 (.PAD(ICACHE_rdata[18]), .C(ICACHE_rdata_i[18]));
		PDIDGZ ipad_ICACHE_rdata19 (.PAD(ICACHE_rdata[19]), .C(ICACHE_rdata_i[19]));
		PDIDGZ ipad_ICACHE_rdata20 (.PAD(ICACHE_rdata[20]), .C(ICACHE_rdata_i[20]));
		PDIDGZ ipad_ICACHE_rdata21 (.PAD(ICACHE_rdata[21]), .C(ICACHE_rdata_i[21]));
		PDIDGZ ipad_ICACHE_rdata22 (.PAD(ICACHE_rdata[22]), .C(ICACHE_rdata_i[22]));
		PDIDGZ ipad_ICACHE_rdata23 (.PAD(ICACHE_rdata[23]), .C(ICACHE_rdata_i[23]));
		PDIDGZ ipad_ICACHE_rdata24 (.PAD(ICACHE_rdata[24]), .C(ICACHE_rdata_i[24]));
		PDIDGZ ipad_ICACHE_rdata25 (.PAD(ICACHE_rdata[25]), .C(ICACHE_rdata_i[25]));
		PDIDGZ ipad_ICACHE_rdata26 (.PAD(ICACHE_rdata[26]), .C(ICACHE_rdata_i[26]));
		PDIDGZ ipad_ICACHE_rdata27 (.PAD(ICACHE_rdata[27]), .C(ICACHE_rdata_i[27]));
		PDIDGZ ipad_ICACHE_rdata28 (.PAD(ICACHE_rdata[28]), .C(ICACHE_rdata_i[28]));
		PDIDGZ ipad_ICACHE_rdata29 (.PAD(ICACHE_rdata[29]), .C(ICACHE_rdata_i[29]));
		PDIDGZ ipad_ICACHE_rdata30 (.PAD(ICACHE_rdata[30]), .C(ICACHE_rdata_i[30]));
		PDIDGZ ipad_ICACHE_rdata31 (.PAD(ICACHE_rdata[31]), .C(ICACHE_rdata_i[31]));
		
		PDIDGZ ipad_DCACHE_rdata0 (.PAD(DCACHE_rdata[0]), .C(DCACHE_rdata_i[0]));
		PDIDGZ ipad_DCACHE_rdata1 (.PAD(DCACHE_rdata[1]), .C(DCACHE_rdata_i[1]));
		PDIDGZ ipad_DCACHE_rdata2 (.PAD(DCACHE_rdata[2]), .C(DCACHE_rdata_i[2]));
		PDIDGZ ipad_DCACHE_rdata3 (.PAD(DCACHE_rdata[3]), .C(DCACHE_rdata_i[3]));
		PDIDGZ ipad_DCACHE_rdata4 (.PAD(DCACHE_rdata[4]), .C(DCACHE_rdata_i[4]));
		PDIDGZ ipad_DCACHE_rdata5 (.PAD(DCACHE_rdata[5]), .C(DCACHE_rdata_i[5]));
		PDIDGZ ipad_DCACHE_rdata6 (.PAD(DCACHE_rdata[6]), .C(DCACHE_rdata_i[6]));
		PDIDGZ ipad_DCACHE_rdata7 (.PAD(DCACHE_rdata[7]), .C(DCACHE_rdata_i[7]));
		PDIDGZ ipad_DCACHE_rdata8 (.PAD(DCACHE_rdata[8]), .C(DCACHE_rdata_i[8]));
		PDIDGZ ipad_DCACHE_rdata9 (.PAD(DCACHE_rdata[9]), .C(DCACHE_rdata_i[9]));
		PDIDGZ ipad_DCACHE_rdata10 (.PAD(DCACHE_rdata[10]), .C(DCACHE_rdata_i[10]));
		PDIDGZ ipad_DCACHE_rdata11 (.PAD(DCACHE_rdata[11]), .C(DCACHE_rdata_i[11]));
		PDIDGZ ipad_DCACHE_rdata12 (.PAD(DCACHE_rdata[12]), .C(DCACHE_rdata_i[12]));
		PDIDGZ ipad_DCACHE_rdata13 (.PAD(DCACHE_rdata[13]), .C(DCACHE_rdata_i[13]));
		PDIDGZ ipad_DCACHE_rdata14 (.PAD(DCACHE_rdata[14]), .C(DCACHE_rdata_i[14]));
		PDIDGZ ipad_DCACHE_rdata15 (.PAD(DCACHE_rdata[15]), .C(DCACHE_rdata_i[15]));
		PDIDGZ ipad_DCACHE_rdata16 (.PAD(DCACHE_rdata[16]), .C(DCACHE_rdata_i[16]));
		PDIDGZ ipad_DCACHE_rdata17 (.PAD(DCACHE_rdata[17]), .C(DCACHE_rdata_i[17]));
		PDIDGZ ipad_DCACHE_rdata18 (.PAD(DCACHE_rdata[18]), .C(DCACHE_rdata_i[18]));
		PDIDGZ ipad_DCACHE_rdata19 (.PAD(DCACHE_rdata[19]), .C(DCACHE_rdata_i[19]));
		PDIDGZ ipad_DCACHE_rdata20 (.PAD(DCACHE_rdata[20]), .C(DCACHE_rdata_i[20]));
		PDIDGZ ipad_DCACHE_rdata21 (.PAD(DCACHE_rdata[21]), .C(DCACHE_rdata_i[21]));
		PDIDGZ ipad_DCACHE_rdata22 (.PAD(DCACHE_rdata[22]), .C(DCACHE_rdata_i[22]));
		PDIDGZ ipad_DCACHE_rdata23 (.PAD(DCACHE_rdata[23]), .C(DCACHE_rdata_i[23]));
		PDIDGZ ipad_DCACHE_rdata24 (.PAD(DCACHE_rdata[24]), .C(DCACHE_rdata_i[24]));
		PDIDGZ ipad_DCACHE_rdata25 (.PAD(DCACHE_rdata[25]), .C(DCACHE_rdata_i[25]));
		PDIDGZ ipad_DCACHE_rdata26 (.PAD(DCACHE_rdata[26]), .C(DCACHE_rdata_i[26]));
		PDIDGZ ipad_DCACHE_rdata27 (.PAD(DCACHE_rdata[27]), .C(DCACHE_rdata_i[27]));
		PDIDGZ ipad_DCACHE_rdata28 (.PAD(DCACHE_rdata[28]), .C(DCACHE_rdata_i[28]));
		PDIDGZ ipad_DCACHE_rdata29 (.PAD(DCACHE_rdata[29]), .C(DCACHE_rdata_i[29]));
		PDIDGZ ipad_DCACHE_rdata30 (.PAD(DCACHE_rdata[30]), .C(DCACHE_rdata_i[30]));
		PDIDGZ ipad_DCACHE_rdata31 (.PAD(DCACHE_rdata[31]), .C(DCACHE_rdata_i[31]));
		
		
		PDO02CDG opad_ICACHE_ren (.PAD(ICACHE_ren), .I(ICACHE_ren_i));
		PDO02CDG opad_ICACHE_wen (.PAD(ICACHE_wen), .I(ICACHE_wen_i));
		PDO02CDG opad_DCACHE_ren (.PAD(DCACHE_ren), .I(DCACHE_ren_i));
		PDO02CDG opad_DCACHE_wen (.PAD(DCACHE_wen), .I(DCACHE_wen_i));
		PDO02CDG opad_test_so (.PAD(test_so), .I(test_so_i));

		PDO02CDG opad_ICACHE_addr0 (.PAD(ICACHE_addr[0]), .I(ICACHE_addr_i[0]));
		PDO02CDG opad_ICACHE_addr1 (.PAD(ICACHE_addr[1]), .I(ICACHE_addr_i[1]));
		PDO02CDG opad_ICACHE_addr2 (.PAD(ICACHE_addr[2]), .I(ICACHE_addr_i[2]));
		PDO02CDG opad_ICACHE_addr3 (.PAD(ICACHE_addr[3]), .I(ICACHE_addr_i[3]));
		PDO02CDG opad_ICACHE_addr4 (.PAD(ICACHE_addr[4]), .I(ICACHE_addr_i[4]));
		PDO02CDG opad_ICACHE_addr5 (.PAD(ICACHE_addr[5]), .I(ICACHE_addr_i[5]));
		PDO02CDG opad_ICACHE_addr6 (.PAD(ICACHE_addr[6]), .I(ICACHE_addr_i[6]));
		PDO02CDG opad_ICACHE_addr7 (.PAD(ICACHE_addr[7]), .I(ICACHE_addr_i[7]));
		PDO02CDG opad_ICACHE_addr8 (.PAD(ICACHE_addr[8]), .I(ICACHE_addr_i[8]));
		PDO02CDG opad_ICACHE_addr9 (.PAD(ICACHE_addr[9]), .I(ICACHE_addr_i[9]));
		PDO02CDG opad_ICACHE_addr10 (.PAD(ICACHE_addr[10]), .I(ICACHE_addr_i[10]));
		PDO02CDG opad_ICACHE_addr11 (.PAD(ICACHE_addr[11]), .I(ICACHE_addr_i[11]));
		PDO02CDG opad_ICACHE_addr12 (.PAD(ICACHE_addr[12]), .I(ICACHE_addr_i[12]));
		PDO02CDG opad_ICACHE_addr13 (.PAD(ICACHE_addr[13]), .I(ICACHE_addr_i[13]));
		PDO02CDG opad_ICACHE_addr14 (.PAD(ICACHE_addr[14]), .I(ICACHE_addr_i[14]));
		PDO02CDG opad_ICACHE_addr15 (.PAD(ICACHE_addr[15]), .I(ICACHE_addr_i[15]));
		PDO02CDG opad_ICACHE_addr16 (.PAD(ICACHE_addr[16]), .I(ICACHE_addr_i[16]));
		PDO02CDG opad_ICACHE_addr17 (.PAD(ICACHE_addr[17]), .I(ICACHE_addr_i[17]));
		PDO02CDG opad_ICACHE_addr18 (.PAD(ICACHE_addr[18]), .I(ICACHE_addr_i[18]));
		PDO02CDG opad_ICACHE_addr19 (.PAD(ICACHE_addr[19]), .I(ICACHE_addr_i[19]));
		PDO02CDG opad_ICACHE_addr20 (.PAD(ICACHE_addr[20]), .I(ICACHE_addr_i[20]));
		PDO02CDG opad_ICACHE_addr21 (.PAD(ICACHE_addr[21]), .I(ICACHE_addr_i[21]));
		PDO02CDG opad_ICACHE_addr22 (.PAD(ICACHE_addr[22]), .I(ICACHE_addr_i[22]));
		PDO02CDG opad_ICACHE_addr23 (.PAD(ICACHE_addr[23]), .I(ICACHE_addr_i[23]));
		PDO02CDG opad_ICACHE_addr24 (.PAD(ICACHE_addr[24]), .I(ICACHE_addr_i[24]));
		PDO02CDG opad_ICACHE_addr25 (.PAD(ICACHE_addr[25]), .I(ICACHE_addr_i[25]));
		PDO02CDG opad_ICACHE_addr26 (.PAD(ICACHE_addr[26]), .I(ICACHE_addr_i[26]));
		PDO02CDG opad_ICACHE_addr27 (.PAD(ICACHE_addr[27]), .I(ICACHE_addr_i[27]));
		PDO02CDG opad_ICACHE_addr28 (.PAD(ICACHE_addr[28]), .I(ICACHE_addr_i[28]));
		PDO02CDG opad_ICACHE_addr29 (.PAD(ICACHE_addr[29]), .I(ICACHE_addr_i[29]));
		PDO02CDG opad_ICACHE_addr30 (.PAD(ICACHE_addr[30]), .I(ICACHE_addr_i[30]));
		PDO02CDG opad_ICACHE_addr31 (.PAD(ICACHE_addr[31]), .I(ICACHE_addr_i[31]));
		
		PDO02CDG opad_DCACHE_addr0 (.PAD(DCACHE_addr[0]), .I(DCACHE_addr_i[0]));
		PDO02CDG opad_DCACHE_addr1 (.PAD(DCACHE_addr[1]), .I(DCACHE_addr_i[1]));
		PDO02CDG opad_DCACHE_addr2 (.PAD(DCACHE_addr[2]), .I(DCACHE_addr_i[2]));
		PDO02CDG opad_DCACHE_addr3 (.PAD(DCACHE_addr[3]), .I(DCACHE_addr_i[3]));
		PDO02CDG opad_DCACHE_addr4 (.PAD(DCACHE_addr[4]), .I(DCACHE_addr_i[4]));
		PDO02CDG opad_DCACHE_addr5 (.PAD(DCACHE_addr[5]), .I(DCACHE_addr_i[5]));
		PDO02CDG opad_DCACHE_addr6 (.PAD(DCACHE_addr[6]), .I(DCACHE_addr_i[6]));
		PDO02CDG opad_DCACHE_addr7 (.PAD(DCACHE_addr[7]), .I(DCACHE_addr_i[7]));
		PDO02CDG opad_DCACHE_addr8 (.PAD(DCACHE_addr[8]), .I(DCACHE_addr_i[8]));
		PDO02CDG opad_DCACHE_addr9 (.PAD(DCACHE_addr[9]), .I(DCACHE_addr_i[9]));
		PDO02CDG opad_DCACHE_addr10 (.PAD(DCACHE_addr[10]), .I(DCACHE_addr_i[10]));
		PDO02CDG opad_DCACHE_addr11 (.PAD(DCACHE_addr[11]), .I(DCACHE_addr_i[11]));
		PDO02CDG opad_DCACHE_addr12 (.PAD(DCACHE_addr[12]), .I(DCACHE_addr_i[12]));
		PDO02CDG opad_DCACHE_addr13 (.PAD(DCACHE_addr[13]), .I(DCACHE_addr_i[13]));
		PDO02CDG opad_DCACHE_addr14 (.PAD(DCACHE_addr[14]), .I(DCACHE_addr_i[14]));
		PDO02CDG opad_DCACHE_addr15 (.PAD(DCACHE_addr[15]), .I(DCACHE_addr_i[15]));
		PDO02CDG opad_DCACHE_addr16 (.PAD(DCACHE_addr[16]), .I(DCACHE_addr_i[16]));
		PDO02CDG opad_DCACHE_addr17 (.PAD(DCACHE_addr[17]), .I(DCACHE_addr_i[17]));
		PDO02CDG opad_DCACHE_addr18 (.PAD(DCACHE_addr[18]), .I(DCACHE_addr_i[18]));
		PDO02CDG opad_DCACHE_addr19 (.PAD(DCACHE_addr[19]), .I(DCACHE_addr_i[19]));
		PDO02CDG opad_DCACHE_addr20 (.PAD(DCACHE_addr[20]), .I(DCACHE_addr_i[20]));
		PDO02CDG opad_DCACHE_addr21 (.PAD(DCACHE_addr[21]), .I(DCACHE_addr_i[21]));
		PDO02CDG opad_DCACHE_addr22 (.PAD(DCACHE_addr[22]), .I(DCACHE_addr_i[22]));
		PDO02CDG opad_DCACHE_addr23 (.PAD(DCACHE_addr[23]), .I(DCACHE_addr_i[23]));
		PDO02CDG opad_DCACHE_addr24 (.PAD(DCACHE_addr[24]), .I(DCACHE_addr_i[24]));
		PDO02CDG opad_DCACHE_addr25 (.PAD(DCACHE_addr[25]), .I(DCACHE_addr_i[25]));
		PDO02CDG opad_DCACHE_addr26 (.PAD(DCACHE_addr[26]), .I(DCACHE_addr_i[26]));
		PDO02CDG opad_DCACHE_addr27 (.PAD(DCACHE_addr[27]), .I(DCACHE_addr_i[27]));
		PDO02CDG opad_DCACHE_addr28 (.PAD(DCACHE_addr[28]), .I(DCACHE_addr_i[28]));
		PDO02CDG opad_DCACHE_addr29 (.PAD(DCACHE_addr[29]), .I(DCACHE_addr_i[29]));
		PDO02CDG opad_DCACHE_addr30 (.PAD(DCACHE_addr[30]), .I(DCACHE_addr_i[30]));
		PDO02CDG opad_DCACHE_addr31 (.PAD(DCACHE_addr[31]), .I(DCACHE_addr_i[31]));
		
		PDO02CDG opad_ICACHE_wdata0 (.PAD(ICACHE_wdata[0]), .I(ICACHE_wdata_i[0]));
		PDO02CDG opad_ICACHE_wdata1 (.PAD(ICACHE_wdata[1]), .I(ICACHE_wdata_i[1]));
		PDO02CDG opad_ICACHE_wdata2 (.PAD(ICACHE_wdata[2]), .I(ICACHE_wdata_i[2]));
		PDO02CDG opad_ICACHE_wdata3 (.PAD(ICACHE_wdata[3]), .I(ICACHE_wdata_i[3]));
		PDO02CDG opad_ICACHE_wdata4 (.PAD(ICACHE_wdata[4]), .I(ICACHE_wdata_i[4]));
		PDO02CDG opad_ICACHE_wdata5 (.PAD(ICACHE_wdata[5]), .I(ICACHE_wdata_i[5]));
		PDO02CDG opad_ICACHE_wdata6 (.PAD(ICACHE_wdata[6]), .I(ICACHE_wdata_i[6]));
		PDO02CDG opad_ICACHE_wdata7 (.PAD(ICACHE_wdata[7]), .I(ICACHE_wdata_i[7]));
		PDO02CDG opad_ICACHE_wdata8 (.PAD(ICACHE_wdata[8]), .I(ICACHE_wdata_i[8]));
		PDO02CDG opad_ICACHE_wdata9 (.PAD(ICACHE_wdata[9]), .I(ICACHE_wdata_i[9]));
		PDO02CDG opad_ICACHE_wdata10 (.PAD(ICACHE_wdata[10]), .I(ICACHE_wdata_i[10]));
		PDO02CDG opad_ICACHE_wdata11 (.PAD(ICACHE_wdata[11]), .I(ICACHE_wdata_i[11]));
		PDO02CDG opad_ICACHE_wdata12 (.PAD(ICACHE_wdata[12]), .I(ICACHE_wdata_i[12]));
		PDO02CDG opad_ICACHE_wdata13 (.PAD(ICACHE_wdata[13]), .I(ICACHE_wdata_i[13]));
		PDO02CDG opad_ICACHE_wdata14 (.PAD(ICACHE_wdata[14]), .I(ICACHE_wdata_i[14]));
		PDO02CDG opad_ICACHE_wdata15 (.PAD(ICACHE_wdata[15]), .I(ICACHE_wdata_i[15]));
		PDO02CDG opad_ICACHE_wdata16 (.PAD(ICACHE_wdata[16]), .I(ICACHE_wdata_i[16]));
		PDO02CDG opad_ICACHE_wdata17 (.PAD(ICACHE_wdata[17]), .I(ICACHE_wdata_i[17]));
		PDO02CDG opad_ICACHE_wdata18 (.PAD(ICACHE_wdata[18]), .I(ICACHE_wdata_i[18]));
		PDO02CDG opad_ICACHE_wdata19 (.PAD(ICACHE_wdata[19]), .I(ICACHE_wdata_i[19]));
		PDO02CDG opad_ICACHE_wdata20 (.PAD(ICACHE_wdata[20]), .I(ICACHE_wdata_i[20]));
		PDO02CDG opad_ICACHE_wdata21 (.PAD(ICACHE_wdata[21]), .I(ICACHE_wdata_i[21]));
		PDO02CDG opad_ICACHE_wdata22 (.PAD(ICACHE_wdata[22]), .I(ICACHE_wdata_i[22]));
		PDO02CDG opad_ICACHE_wdata23 (.PAD(ICACHE_wdata[23]), .I(ICACHE_wdata_i[23]));
		PDO02CDG opad_ICACHE_wdata24 (.PAD(ICACHE_wdata[24]), .I(ICACHE_wdata_i[24]));
		PDO02CDG opad_ICACHE_wdata25 (.PAD(ICACHE_wdata[25]), .I(ICACHE_wdata_i[25]));
		PDO02CDG opad_ICACHE_wdata26 (.PAD(ICACHE_wdata[26]), .I(ICACHE_wdata_i[26]));
		PDO02CDG opad_ICACHE_wdata27 (.PAD(ICACHE_wdata[27]), .I(ICACHE_wdata_i[27]));
		PDO02CDG opad_ICACHE_wdata28 (.PAD(ICACHE_wdata[28]), .I(ICACHE_wdata_i[28]));
		PDO02CDG opad_ICACHE_wdata29 (.PAD(ICACHE_wdata[29]), .I(ICACHE_wdata_i[29]));
		PDO02CDG opad_ICACHE_wdata30 (.PAD(ICACHE_wdata[30]), .I(ICACHE_wdata_i[30]));
		PDO02CDG opad_ICACHE_wdata31 (.PAD(ICACHE_wdata[31]), .I(ICACHE_wdata_i[31]));
		
		PDO02CDG opad_DCACHE_wdata0 (.PAD(DCACHE_wdata[0]), .I(DCACHE_wdata_i[0]));
		PDO02CDG opad_DCACHE_wdata1 (.PAD(DCACHE_wdata[1]), .I(DCACHE_wdata_i[1]));
		PDO02CDG opad_DCACHE_wdata2 (.PAD(DCACHE_wdata[2]), .I(DCACHE_wdata_i[2]));
		PDO02CDG opad_DCACHE_wdata3 (.PAD(DCACHE_wdata[3]), .I(DCACHE_wdata_i[3]));
		PDO02CDG opad_DCACHE_wdata4 (.PAD(DCACHE_wdata[4]), .I(DCACHE_wdata_i[4]));
		PDO02CDG opad_DCACHE_wdata5 (.PAD(DCACHE_wdata[5]), .I(DCACHE_wdata_i[5]));
		PDO02CDG opad_DCACHE_wdata6 (.PAD(DCACHE_wdata[6]), .I(DCACHE_wdata_i[6]));
		PDO02CDG opad_DCACHE_wdata7 (.PAD(DCACHE_wdata[7]), .I(DCACHE_wdata_i[7]));
		PDO02CDG opad_DCACHE_wdata8 (.PAD(DCACHE_wdata[8]), .I(DCACHE_wdata_i[8]));
		PDO02CDG opad_DCACHE_wdata9 (.PAD(DCACHE_wdata[9]), .I(DCACHE_wdata_i[9]));
		PDO02CDG opad_DCACHE_wdata10 (.PAD(DCACHE_wdata[10]), .I(DCACHE_wdata_i[10]));
		PDO02CDG opad_DCACHE_wdata11 (.PAD(DCACHE_wdata[11]), .I(DCACHE_wdata_i[11]));
		PDO02CDG opad_DCACHE_wdata12 (.PAD(DCACHE_wdata[12]), .I(DCACHE_wdata_i[12]));
		PDO02CDG opad_DCACHE_wdata13 (.PAD(DCACHE_wdata[13]), .I(DCACHE_wdata_i[13]));
		PDO02CDG opad_DCACHE_wdata14 (.PAD(DCACHE_wdata[14]), .I(DCACHE_wdata_i[14]));
		PDO02CDG opad_DCACHE_wdata15 (.PAD(DCACHE_wdata[15]), .I(DCACHE_wdata_i[15]));
		PDO02CDG opad_DCACHE_wdata16 (.PAD(DCACHE_wdata[16]), .I(DCACHE_wdata_i[16]));
		PDO02CDG opad_DCACHE_wdata17 (.PAD(DCACHE_wdata[17]), .I(DCACHE_wdata_i[17]));
		PDO02CDG opad_DCACHE_wdata18 (.PAD(DCACHE_wdata[18]), .I(DCACHE_wdata_i[18]));
		PDO02CDG opad_DCACHE_wdata19 (.PAD(DCACHE_wdata[19]), .I(DCACHE_wdata_i[19]));
		PDO02CDG opad_DCACHE_wdata20 (.PAD(DCACHE_wdata[20]), .I(DCACHE_wdata_i[20]));
		PDO02CDG opad_DCACHE_wdata21 (.PAD(DCACHE_wdata[21]), .I(DCACHE_wdata_i[21]));
		PDO02CDG opad_DCACHE_wdata22 (.PAD(DCACHE_wdata[22]), .I(DCACHE_wdata_i[22]));
		PDO02CDG opad_DCACHE_wdata23 (.PAD(DCACHE_wdata[23]), .I(DCACHE_wdata_i[23]));
		PDO02CDG opad_DCACHE_wdata24 (.PAD(DCACHE_wdata[24]), .I(DCACHE_wdata_i[24]));
		PDO02CDG opad_DCACHE_wdata25 (.PAD(DCACHE_wdata[25]), .I(DCACHE_wdata_i[25]));
		PDO02CDG opad_DCACHE_wdata26 (.PAD(DCACHE_wdata[26]), .I(DCACHE_wdata_i[26]));
		PDO02CDG opad_DCACHE_wdata27 (.PAD(DCACHE_wdata[27]), .I(DCACHE_wdata_i[27]));
		PDO02CDG opad_DCACHE_wdata28 (.PAD(DCACHE_wdata[28]), .I(DCACHE_wdata_i[28]));
		PDO02CDG opad_DCACHE_wdata29 (.PAD(DCACHE_wdata[29]), .I(DCACHE_wdata_i[29]));
		PDO02CDG opad_DCACHE_wdata30 (.PAD(DCACHE_wdata[30]), .I(DCACHE_wdata_i[30]));
		PDO02CDG opad_DCACHE_wdata31 (.PAD(DCACHE_wdata[31]), .I(DCACHE_wdata_i[31]));
		
		MIPS_Pipeline MIPS( clk_i, rst_i, ICACHE_addr_i, ICACHE_rdata_i, ICACHE_ren_i, 
							ICACHE_wen_i, ICACHE_wdata_i, ICACHE_stall_i, DCACHE_addr_i, DCACHE_rdata_i, 
							DCACHE_ren_i, DCACHE_wen_i, DCACHE_wdata_i, DCACHE_stall_i, test_si_i, test_so_i, 
							test_se_i );
		
endmodule 