* SPICE NETLIST
***************************************

.SUBCKT NC1 ng nds
.ENDS
***************************************
.SUBCKT NC2 ng nds
.ENDS
***************************************
.SUBCKT PC1 ng nds
.ENDS
***************************************
.SUBCKT PC2 ng nds
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_2
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_3
** N=10 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_4
** N=11 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_5
** N=12 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_6
** N=21 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_7
** N=19 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_8
** N=18 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_9
** N=17 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_10
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_11
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_12
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_13
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT PDIDGZ C PAD
** N=3 EP=2 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_14 1 2 3 4 5 6 7 8 9 10 13
** N=13 EP=11 IP=15 FDC=0
X0 1 6 PDIDGZ $T=2600000 2155570 0 90 $X=2354000 $Y=2160848
X1 2 7 PDIDGZ $T=2600000 2195255 0 90 $X=2354000 $Y=2200533
X2 3 8 PDIDGZ $T=2600000 2234940 0 90 $X=2354000 $Y=2240218
X3 4 9 PDIDGZ $T=2600000 2274625 0 90 $X=2354000 $Y=2279903
X4 5 10 PDIDGZ $T=2600000 2314310 0 90 $X=2354000 $Y=2319588
.ENDS
***************************************
.SUBCKT ICV_15 1 2 3 4 5 6 7 8 9 10 15
** N=15 EP=11 IP=15 FDC=0
X0 1 6 PDIDGZ $T=2600000 1957145 0 90 $X=2354000 $Y=1962423
X1 2 7 PDIDGZ $T=2600000 1996830 0 90 $X=2354000 $Y=2002108
X2 3 8 PDIDGZ $T=2600000 2036515 0 90 $X=2354000 $Y=2041793
X3 4 9 PDIDGZ $T=2600000 2076200 0 90 $X=2354000 $Y=2081478
X4 5 10 PDIDGZ $T=2600000 2115885 0 90 $X=2354000 $Y=2121163
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3 4 5 6 7 8 9 10 13
** N=13 EP=11 IP=15 FDC=0
X0 1 6 PDIDGZ $T=2600000 1758720 0 90 $X=2354000 $Y=1763998
X1 2 7 PDIDGZ $T=2600000 1798405 0 90 $X=2354000 $Y=1803683
X2 3 8 PDIDGZ $T=2600000 1838090 0 90 $X=2354000 $Y=1843368
X3 4 9 PDIDGZ $T=2600000 1877775 0 90 $X=2354000 $Y=1883053
X4 5 10 PDIDGZ $T=2600000 1917460 0 90 $X=2354000 $Y=1922738
.ENDS
***************************************
.SUBCKT PDO02CDG I PAD
** N=3 EP=2 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_17 1 2 3 4 5 6 7 8 9 12 13 14 15 16 17 18 19 20 29
** N=30 EP=19 IP=27 FDC=0
X0 3 17 PDIDGZ $T=2600000 1599980 0 90 $X=2354000 $Y=1605258
X1 4 18 PDIDGZ $T=2600000 1639665 0 90 $X=2354000 $Y=1644943
X2 5 19 PDIDGZ $T=2600000 1679350 0 90 $X=2354000 $Y=1684628
X3 2 20 PDIDGZ $T=2600000 1719035 0 90 $X=2354000 $Y=1724313
X4 6 12 PDO02CDG $T=2600000 1401555 0 90 $X=2354000 $Y=1405243
X5 7 13 PDO02CDG $T=2600000 1441240 0 90 $X=2354000 $Y=1444928
X6 1 14 PDO02CDG $T=2600000 1480925 0 90 $X=2354000 $Y=1484613
X7 8 15 PDO02CDG $T=2600000 1520610 0 90 $X=2354000 $Y=1524298
X8 9 16 PDO02CDG $T=2600000 1560295 0 90 $X=2354000 $Y=1563983
.ENDS
***************************************
.SUBCKT ICV_18 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 24
** N=24 EP=17 IP=24 FDC=0
X0 1 9 PDO02CDG $T=2600000 1004705 0 90 $X=2354000 $Y=1008393
X1 2 10 PDO02CDG $T=2600000 1044390 0 90 $X=2354000 $Y=1048078
X2 3 11 PDO02CDG $T=2600000 1084075 0 90 $X=2354000 $Y=1087763
X3 4 12 PDO02CDG $T=2600000 1123760 0 90 $X=2354000 $Y=1127448
X4 5 13 PDO02CDG $T=2600000 1163445 0 90 $X=2354000 $Y=1167133
X5 6 14 PDO02CDG $T=2600000 1203130 0 90 $X=2354000 $Y=1206818
X6 7 15 PDO02CDG $T=2600000 1242815 0 90 $X=2354000 $Y=1246503
X7 8 16 PDO02CDG $T=2600000 1282500 0 90 $X=2354000 $Y=1286188
.ENDS
***************************************
.SUBCKT ICV_19 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 23
** N=23 EP=19 IP=27 FDC=0
X0 2 10 PDO02CDG $T=2600000 647540 0 90 $X=2354000 $Y=651228
X1 3 11 PDO02CDG $T=2600000 687225 0 90 $X=2354000 $Y=690913
X2 4 12 PDO02CDG $T=2600000 726910 0 90 $X=2354000 $Y=730598
X3 1 13 PDO02CDG $T=2600000 766595 0 90 $X=2354000 $Y=770283
X4 5 14 PDO02CDG $T=2600000 806280 0 90 $X=2354000 $Y=809968
X5 6 15 PDO02CDG $T=2600000 845965 0 90 $X=2354000 $Y=849653
X6 7 16 PDO02CDG $T=2600000 885650 0 90 $X=2354000 $Y=889338
X7 8 17 PDO02CDG $T=2600000 925335 0 90 $X=2354000 $Y=929023
X8 9 18 PDO02CDG $T=2600000 965020 0 90 $X=2354000 $Y=968708
.ENDS
***************************************
.SUBCKT ICV_20 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 26
** N=26 EP=21 IP=30 FDC=0
X0 1 11 PDO02CDG $T=2600000 250690 0 90 $X=2354000 $Y=254378
X1 2 12 PDO02CDG $T=2600000 290375 0 90 $X=2354000 $Y=294063
X2 3 13 PDO02CDG $T=2600000 330060 0 90 $X=2354000 $Y=333748
X3 4 14 PDO02CDG $T=2600000 369745 0 90 $X=2354000 $Y=373433
X4 5 15 PDO02CDG $T=2600000 409430 0 90 $X=2354000 $Y=413118
X5 6 16 PDO02CDG $T=2600000 449115 0 90 $X=2354000 $Y=452803
X6 7 17 PDO02CDG $T=2600000 488800 0 90 $X=2354000 $Y=492488
X7 8 18 PDO02CDG $T=2600000 528485 0 90 $X=2354000 $Y=532173
X8 9 19 PDO02CDG $T=2600000 568170 0 90 $X=2354000 $Y=571858
X9 10 20 PDO02CDG $T=2600000 607855 0 90 $X=2354000 $Y=611543
.ENDS
***************************************
.SUBCKT ICV_21
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_22
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_23
** N=82 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_24 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 81 82 83 84
+ 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104
+ 105 106 135
** N=135 EP=103 IP=153 FDC=0
X0 1 52 PDIDGZ $T=285690 2600000 0 180 $X=255970 $Y=2354000
X1 2 53 PDIDGZ $T=325375 2600000 0 180 $X=295655 $Y=2354000
X2 3 54 PDIDGZ $T=365060 2600000 0 180 $X=335340 $Y=2354000
X3 4 55 PDIDGZ $T=404745 2600000 0 180 $X=375025 $Y=2354000
X4 5 56 PDIDGZ $T=444430 2600000 0 180 $X=414710 $Y=2354000
X5 6 57 PDIDGZ $T=484115 2600000 0 180 $X=454395 $Y=2354000
X6 7 58 PDIDGZ $T=523800 2600000 0 180 $X=494080 $Y=2354000
X7 8 59 PDIDGZ $T=563485 2600000 0 180 $X=533765 $Y=2354000
X8 9 60 PDIDGZ $T=603170 2600000 0 180 $X=573450 $Y=2354000
X9 10 61 PDIDGZ $T=642855 2600000 0 180 $X=613135 $Y=2354000
X10 11 62 PDIDGZ $T=682540 2600000 0 180 $X=652820 $Y=2354000
X11 12 63 PDIDGZ $T=722225 2600000 0 180 $X=692505 $Y=2354000
X12 13 64 PDIDGZ $T=761910 2600000 0 180 $X=732190 $Y=2354000
X13 14 65 PDIDGZ $T=801595 2600000 0 180 $X=771875 $Y=2354000
X14 15 66 PDIDGZ $T=841280 2600000 0 180 $X=811560 $Y=2354000
X15 16 67 PDIDGZ $T=880965 2600000 0 180 $X=851245 $Y=2354000
X16 17 68 PDIDGZ $T=920650 2600000 0 180 $X=890930 $Y=2354000
X17 18 69 PDIDGZ $T=960335 2600000 0 180 $X=930615 $Y=2354000
X18 19 70 PDIDGZ $T=1000020 2600000 0 180 $X=970300 $Y=2354000
X19 20 71 PDIDGZ $T=1039705 2600000 0 180 $X=1009985 $Y=2354000
X20 21 72 PDIDGZ $T=1079390 2600000 0 180 $X=1049670 $Y=2354000
X21 22 73 PDIDGZ $T=1119075 2600000 0 180 $X=1089355 $Y=2354000
X22 23 74 PDIDGZ $T=1158760 2600000 0 180 $X=1129040 $Y=2354000
X23 24 75 PDIDGZ $T=1198445 2600000 0 180 $X=1168725 $Y=2354000
X24 25 76 PDIDGZ $T=1238130 2600000 0 180 $X=1208410 $Y=2354000
X25 26 81 PDIDGZ $T=1357185 2600000 0 180 $X=1327465 $Y=2354000
X26 27 82 PDIDGZ $T=1396870 2600000 0 180 $X=1367150 $Y=2354000
X27 28 83 PDIDGZ $T=1436555 2600000 0 180 $X=1406835 $Y=2354000
X28 29 84 PDIDGZ $T=1476240 2600000 0 180 $X=1446520 $Y=2354000
X29 30 85 PDIDGZ $T=1515925 2600000 0 180 $X=1486205 $Y=2354000
X30 31 86 PDIDGZ $T=1555610 2600000 0 180 $X=1525890 $Y=2354000
X31 32 87 PDIDGZ $T=1595295 2600000 0 180 $X=1565575 $Y=2354000
X32 33 88 PDIDGZ $T=1634980 2600000 0 180 $X=1605260 $Y=2354000
X33 34 89 PDIDGZ $T=1674665 2600000 0 180 $X=1644945 $Y=2354000
X34 35 90 PDIDGZ $T=1714350 2600000 0 180 $X=1684630 $Y=2354000
X35 36 91 PDIDGZ $T=1754035 2600000 0 180 $X=1724315 $Y=2354000
X36 37 92 PDIDGZ $T=1793720 2600000 0 180 $X=1764000 $Y=2354000
X37 38 93 PDIDGZ $T=1833405 2600000 0 180 $X=1803685 $Y=2354000
X38 39 94 PDIDGZ $T=1873090 2600000 0 180 $X=1843370 $Y=2354000
X39 40 95 PDIDGZ $T=1912775 2600000 0 180 $X=1883055 $Y=2354000
X40 41 96 PDIDGZ $T=1952460 2600000 0 180 $X=1922740 $Y=2354000
X41 42 97 PDIDGZ $T=1992145 2600000 0 180 $X=1962425 $Y=2354000
X42 43 98 PDIDGZ $T=2031830 2600000 0 180 $X=2002110 $Y=2354000
X43 44 99 PDIDGZ $T=2071515 2600000 0 180 $X=2041795 $Y=2354000
X44 45 100 PDIDGZ $T=2111200 2600000 0 180 $X=2081480 $Y=2354000
X45 46 101 PDIDGZ $T=2150885 2600000 0 180 $X=2121165 $Y=2354000
X46 47 102 PDIDGZ $T=2190570 2600000 0 180 $X=2160850 $Y=2354000
X47 48 103 PDIDGZ $T=2230255 2600000 0 180 $X=2200535 $Y=2354000
X48 49 104 PDIDGZ $T=2269940 2600000 0 180 $X=2240220 $Y=2354000
X49 50 105 PDIDGZ $T=2309625 2600000 0 180 $X=2279905 $Y=2354000
X50 51 106 PDIDGZ $T=2349310 2600000 0 180 $X=2319590 $Y=2354000
.ENDS
***************************************
.SUBCKT ICV_25
** N=75902 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_26
** N=72534 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR2X1 A B VSS VDD Y
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT TIELO VDD VSS Y
** N=4 EP=3 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKINVX20 A VSS Y VDD
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_27 28 29 63 64 66 168 169 184 187 188 4159
** N=90492 EP=11 IP=23 FDC=0
X0 188 187 28 29 184 OR2X1 $T=1705220 1849510 0 180 $X=1703380 $Y=1845570
X1 29 28 63 TIELO $T=746120 1849510 0 0 $X=746118 $Y=1849258
X2 29 28 64 TIELO $T=747040 1849510 0 0 $X=747038 $Y=1849258
X3 29 28 66 TIELO $T=747960 1849510 0 0 $X=747958 $Y=1849258
X4 169 28 168 29 CLKINVX20 $T=1571820 1849510 0 0 $X=1571818 $Y=1849258
.ENDS
***************************************
.SUBCKT TIEHI VDD VSS Y
** N=4 EP=3 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUFX12 A Y VSS VDD
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR2BX1 AN B VDD VSS Y
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKBUFX3 A VSS Y VDD
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI2BB2XL A0N A1N B1 VSS B0 VDD Y
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKBUFX4 A Y VSS VDD
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT SDFFRXL SE D SI CK RN QN VDD VSS Q
** N=10 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKBUFX2 A VSS Y VDD
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MX2XL S0 B A VSS VDD Y
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MXI2X1 B S0 Y A VSS VDD
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AND2X2 A VDD B VSS Y
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AND2XL A B VSS VDD Y
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND2X1 B VSS A Y VDD
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT SDFFNSRXL SE SI D CKN RN SN QN VSS VDD Q
** N=11 EP=10 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR2X1 B VDD A Y VSS
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKINVX1 A VSS VDD Y
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INVXL A VDD VSS Y
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INVX1 A VSS VDD Y
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKINVX3 A VSS Y VDD
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ANTENNA VSS VDD A
** N=4 EP=3 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKBUFX20 A VSS Y VDD
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_28 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15
** N=15 EP=15 IP=18 FDC=0
X0 3 2 4 5 6 1 MXI2X1 $T=0 0 0 0 $X=-2 $Y=-252
X1 7 8 9 10 11 12 13 6 1 14 SDFFNSRXL $T=3220 0 0 0 $X=3218 $Y=-252
.ENDS
***************************************
.SUBCKT MXI4X1 A B S0 D C S1 VSS Y VDD
** N=10 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKINVX12 A VSS Y VDD
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MXI4XL A B S0 D C S1 VSS Y VDD
** N=10 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_29 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15
** N=15 EP=15 IP=18 FDC=0
X0 3 2 4 5 6 1 MXI2X1 $T=0 0 0 0 $X=-2 $Y=-252
X1 7 8 9 10 11 12 13 6 1 14 SDFFNSRXL $T=4140 0 0 0 $X=4138 $Y=-252
.ENDS
***************************************
.SUBCKT MX4X1 C D S0 B A S1 VDD VSS Y
** N=10 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MXI2X2 S0 B Y A VSS VDD
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INVX12 A Y VDD VSS
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKMX2X2 S0 B A VDD VSS Y
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INVX2 A VSS VDD Y
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKINVX8 A VSS Y VDD
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MX4XL C D S0 B A S1 VDD VSS Y
** N=10 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR2XL B VDD A Y VSS
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR2BXL AN B VDD VSS Y
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INVX3 A Y VSS VDD
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKBUFX16 A VSS Y VDD
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND2XL B VSS A Y VDD
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI221XL B1 B0 VSS A0 A1 VDD C0 Y
** N=9 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OA22X1 A1 A0 B0 B1 VSS VDD Y
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AO22X1 B1 B0 A0 VSS A1 VDD Y
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR4X1 D VDD C B A VSS Y
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND3BX1 AN VDD VSS C B Y
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XOR2X1 A B Y VSS VDD
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI21XL A1 A0 VSS B0 VDD Y
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MX2X1 S0 B A VSS VDD Y
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XOR2XL A B Y VSS VDD
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI222XL C0 C1 VDD B1 B0 A0 A1 Y VSS
** N=10 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AO21X1 A1 A0 B0 VSS VDD Y
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI22XL B1 B0 VDD A0 A1 VSS Y
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XOR3X1 A B C VDD Y VSS
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND2BXL AN B VSS VDD Y
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ADDFXL B A CI CO VDD VSS S
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT SDFFRX2 D SE SI CK RN QN Q VDD VSS
** N=10 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI211X1 A1 A0 VSS C0 VDD B0 Y
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI2BB2X1 A1N A0N B1 VDD B0 Y VSS
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XNOR2X1 A B Y VDD VSS
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR3X1 C VDD B VSS A Y
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AND4X1 A B C VSS D VDD Y
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AO21XL A1 A0 B0 VSS VDD Y
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI21X1 A1 A0 VDD B0 VSS Y
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI22X1 B1 B0 VDD A0 A1 VSS Y
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND2BX1 AN B VSS Y VDD
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OA21XL A1 A0 B0 VSS VDD Y
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XNOR2XL A B Y VSS VDD
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI31XL VSS A2 A1 A0 B0 Y VDD
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CMPR32X2 B A C CO VSS VDD S
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND3BXL AN C VSS B VDD Y
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI2BB1X1 A0N A1N B0 VDD VSS Y
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT SDFFRHQX8 CK SE D SI RN Q VSS VDD
** N=9 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND4BBXL BN D C Y VDD AN VSS
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUFX2 A Y VSS VDD
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND4XL D VSS C B A Y VDD
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT SDFFSXL SE SI D CK SN QN VSS VDD Q
** N=10 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT TLATX1 G D Q VDD VSS QN
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT SDFFRX4 D SE SI CK RN QN Q VDD VSS
** N=10 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI22XL B1 VSS B0 A0 A1 Y VDD
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AND3XL A B VSS C VDD Y
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND3XL C VSS B VDD A Y
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI32X1 A2 A1 VSS A0 B0 Y VDD B1
** N=9 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI2BB1X1 A1N A0N B0 VSS Y VDD
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR3XL C VDD B VSS A Y
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AO22XL B1 B0 A0 A1 VSS VDD Y
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND3X1 C VSS B VDD A Y
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR4XL D VDD C B Y VSS A
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND4X1 D VSS C B A Y VDD
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI2BB2XL A1N A0N VDD B1 B0 VSS Y
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR4BX1 AN D VDD C B Y VSS
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AND3X2 A B C VSS VDD Y
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI211X1 A1 VDD A0 C0 VSS B0 Y
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND4BX1 AN D VSS C B Y VDD
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR3XL A B C VDD VSS Y
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR4X1 A B C D VDD VSS Y
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR3X2 A B C VDD VSS Y
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI211XL A1 VDD A0 C0 VSS B0 Y
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI221XL B1 B0 VDD A0 A1 VSS C0 Y
** N=9 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUFX4 A VSS VDD Y
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI33X1 B2 B1 B0 VSS A0 A1 A2 VDD Y
** N=10 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI2BB1XL A1N A0N B0 VSS VDD Y
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKBUFX8 A VSS Y VDD
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_30 2 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202
+ 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242
+ 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261 262
+ 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281 282
+ 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300 301 302
+ 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322
+ 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342
+ 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362
+ 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382
+ 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402
+ 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422
+ 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442
+ 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462
+ 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482
+ 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502
+ 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522
+ 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542
+ 543 544 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562
+ 563 564 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582
+ 583 584 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602
+ 603 604 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622
+ 623 624 625 626 627 628 629 630 631 3961
** N=193159 EP=610 IP=22561 FDC=0
X0 10280 10169 24 25 10275 OR2X1 $T=1139880 1495270 0 180 $X=1138040 $Y=1491330
X1 10387 10599 24 25 10594 OR2X1 $T=1165180 1510030 0 180 $X=1163340 $Y=1506090
X2 10817 11179 24 25 11184 OR2X1 $T=1201980 1465750 0 0 $X=1201978 $Y=1465498
X3 11312 193 24 25 11374 OR2X1 $T=1213480 1355050 1 0 $X=1213478 $Y=1351110
X4 11526 11475 24 25 11232 OR2X1 $T=1227280 1391950 0 180 $X=1225440 $Y=1388010
X5 11455 11387 24 25 11501 OR2X1 $T=1225900 1399330 0 0 $X=1225898 $Y=1399078
X6 10644 11498 24 25 11508 OR2X1 $T=1226360 1369810 1 0 $X=1226358 $Y=1365870
X7 11581 11588 24 25 11651 OR2X1 $T=1231880 1362430 1 0 $X=1231878 $Y=1358490
X8 11018 92 24 25 11617 OR2X1 $T=1232800 1458370 0 0 $X=1232798 $Y=1458118
X9 219 220 24 25 11754 OR2X1 $T=1243840 1355050 1 0 $X=1243838 $Y=1351110
X10 11872 11812 24 25 11756 OR2X1 $T=1249820 1473130 1 180 $X=1247980 $Y=1472878
X11 15168 15158 24 25 15152 OR2X1 $T=1556640 1450990 1 180 $X=1554800 $Y=1450738
X12 25 24 2 TIELO $T=746120 1731430 1 0 $X=746118 $Y=1727490
X13 25 24 630 TIELO $T=1852880 1524790 0 0 $X=1852878 $Y=1524538
X14 25 24 12615 TIEHI $T=1343660 1473130 0 0 $X=1343658 $Y=1472878
X15 25 24 12342 TIEHI $T=1376780 1532170 1 0 $X=1376778 $Y=1528230
X16 25 24 12507 TIEHI $T=1380000 1384570 0 0 $X=1379998 $Y=1384318
X17 25 24 13267 TIEHI $T=1380460 1569070 1 0 $X=1380458 $Y=1565130
X18 25 24 12399 TIEHI $T=1381840 1473130 1 0 $X=1381838 $Y=1469190
X19 25 24 12721 TIEHI $T=1381840 1517410 1 0 $X=1381838 $Y=1513470
X20 25 24 12506 TIEHI $T=1384600 1369810 0 0 $X=1384598 $Y=1369558
X21 25 24 12462 TIEHI $T=1385060 1406710 0 0 $X=1385058 $Y=1406458
X22 25 24 12497 TIEHI $T=1385060 1539550 1 0 $X=1385058 $Y=1535610
X23 25 24 12398 TIEHI $T=1386900 1428850 1 0 $X=1386898 $Y=1424910
X24 25 24 12508 TIEHI $T=1389660 1450990 1 0 $X=1389658 $Y=1447050
X25 25 24 12560 TIEHI $T=1391960 1458370 0 0 $X=1391958 $Y=1458118
X26 25 24 12688 TIEHI $T=1395640 1436230 0 0 $X=1395638 $Y=1435978
X27 25 24 12805 TIEHI $T=1396560 1554310 0 0 $X=1396558 $Y=1554058
X28 25 24 12684 TIEHI $T=1403000 1502650 0 0 $X=1402998 $Y=1502398
X29 25 24 12683 TIEHI $T=1405760 1377190 0 0 $X=1405758 $Y=1376938
X30 25 24 12687 TIEHI $T=1405760 1414090 0 0 $X=1405758 $Y=1413838
X31 25 24 12692 TIEHI $T=1409440 1546930 0 0 $X=1409438 $Y=1546678
X32 25 24 12818 TIEHI $T=1413580 1362430 1 0 $X=1413578 $Y=1358490
X33 25 24 12678 TIEHI $T=1414960 1487890 0 0 $X=1414958 $Y=1487638
X34 25 24 12679 TIEHI $T=1418640 1495270 0 0 $X=1418638 $Y=1495018
X35 25 24 12787 TIEHI $T=1420020 1443610 0 0 $X=1420018 $Y=1443358
X36 25 24 12926 TIEHI $T=1425540 1399330 1 0 $X=1425538 $Y=1395390
X37 25 24 12974 TIEHI $T=1430600 1546930 0 0 $X=1430598 $Y=1546678
X38 25 24 12925 TIEHI $T=1431060 1465750 0 0 $X=1431058 $Y=1465498
X39 25 24 13025 TIEHI $T=1436580 1510030 1 0 $X=1436578 $Y=1506090
X40 25 24 13042 TIEHI $T=1437040 1524790 0 0 $X=1437038 $Y=1524538
X41 25 24 13062 TIEHI $T=1437500 1532170 0 0 $X=1437498 $Y=1531918
X42 25 24 13096 TIEHI $T=1443480 1517410 1 0 $X=1443478 $Y=1513470
X43 25 24 13152 TIEHI $T=1450380 1436230 0 0 $X=1450378 $Y=1435978
X44 25 24 13391 TIEHI $T=1464180 1406710 1 0 $X=1464178 $Y=1402770
X45 25 24 13383 TIEHI $T=1465100 1428850 1 0 $X=1465098 $Y=1424910
X46 25 24 13397 TIEHI $T=1465100 1495270 1 0 $X=1465098 $Y=1491330
X47 25 24 13413 TIEHI $T=1465560 1495270 0 0 $X=1465558 $Y=1495018
X48 25 24 13425 TIEHI $T=1475220 1473130 0 0 $X=1475218 $Y=1472878
X49 25 24 441 TIEHI $T=1477520 1355050 1 0 $X=1477518 $Y=1351110
X50 25 24 13475 TIEHI $T=1478440 1362430 1 0 $X=1478438 $Y=1358490
X51 25 24 13530 TIEHI $T=1478440 1414090 1 0 $X=1478438 $Y=1410150
X52 25 24 13476 TIEHI $T=1478900 1384570 1 0 $X=1478898 $Y=1380630
X53 25 24 13485 TIEHI $T=1479360 1391950 1 0 $X=1479358 $Y=1388010
X54 25 24 13576 TIEHI $T=1481660 1458370 1 0 $X=1481658 $Y=1454430
X55 25 24 13503 TIEHI $T=1486720 1421470 1 0 $X=1486718 $Y=1417530
X56 25 24 13655 TIEHI $T=1487180 1377190 1 0 $X=1487178 $Y=1373250
X57 25 24 13651 TIEHI $T=1488560 1480510 0 0 $X=1488558 $Y=1480258
X58 25 24 13668 TIEHI $T=1489480 1450990 1 0 $X=1489478 $Y=1447050
X59 25 24 631 TIEHI $T=1852880 1561690 0 0 $X=1852878 $Y=1561438
X60 16194 628 24 25 BUFX12 $T=1840000 1443610 1 0 $X=1839998 $Y=1439670
X61 16091 629 24 25 BUFX12 $T=1841840 1458370 1 0 $X=1841838 $Y=1454430
X62 35 9745 25 24 9739 NOR2BX1 $T=1106760 1391950 0 180 $X=1104920 $Y=1388010
X63 10490 10460 25 24 10274 NOR2BX1 $T=1152300 1495270 0 180 $X=1150460 $Y=1491330
X64 10455 10389 25 24 119 NOR2BX1 $T=1153680 1473130 1 0 $X=1153678 $Y=1469190
X65 11541 92 25 24 11626 NOR2BX1 $T=1233720 1458370 1 0 $X=1233718 $Y=1454430
X66 11313 11469 25 24 11660 NOR2BX1 $T=1234180 1414090 1 0 $X=1234178 $Y=1410150
X67 11692 12206 25 24 12179 NOR2BX1 $T=1275120 1487890 0 180 $X=1273280 $Y=1483950
X68 76 10937 25 24 12670 NOR2BX1 $T=1302720 1362430 0 0 $X=1302718 $Y=1362178
X69 10033 10137 25 24 12693 NOR2BX1 $T=1311460 1355050 0 0 $X=1311458 $Y=1354798
X70 10137 10033 25 24 12778 NOR2BX1 $T=1318820 1362430 1 0 $X=1318818 $Y=1358490
X71 386 14915 25 24 14854 NOR2BX1 $T=1530880 1443610 0 180 $X=1529040 $Y=1439670
X72 537 550 25 24 14937 NOR2BX1 $T=1537780 1355050 0 180 $X=1535940 $Y=1351110
X73 537 14915 25 24 14882 NOR2BX1 $T=1538700 1443610 1 180 $X=1536860 $Y=1443358
X74 391 14969 25 24 14957 NOR2BX1 $T=1538700 1458370 1 180 $X=1536860 $Y=1458118
X75 360 14981 25 24 14941 NOR2BX1 $T=1540080 1450990 1 180 $X=1538240 $Y=1450738
X76 339 15066 25 24 14960 NOR2BX1 $T=1544220 1377190 1 180 $X=1542380 $Y=1376938
X77 382 15066 25 24 15067 NOR2BX1 $T=1548820 1377190 1 180 $X=1546980 $Y=1376938
X78 537 14981 25 24 15091 NOR2BX1 $T=1551120 1458370 0 180 $X=1549280 $Y=1454430
X79 339 14989 25 24 15061 NOR2BX1 $T=1551580 1414090 0 180 $X=1549740 $Y=1410150
X80 374 14989 25 24 15062 NOR2BX1 $T=1551580 1414090 1 180 $X=1549740 $Y=1413838
X81 339 14969 25 24 15129 NOR2BX1 $T=1552960 1465750 0 180 $X=1551120 $Y=1461810
X82 357 15185 25 24 15175 NOR2BX1 $T=1559400 1406710 1 0 $X=1559398 $Y=1402770
X83 15243 386 25 24 15159 NOR2BX1 $T=1561240 1377190 0 180 $X=1559400 $Y=1373250
X84 401 15280 25 24 15236 NOR2BX1 $T=1564000 1458370 0 180 $X=1562160 $Y=1454430
X85 537 15185 25 24 15238 NOR2BX1 $T=1565840 1406710 1 180 $X=1564000 $Y=1406458
X86 401 15266 25 24 15263 NOR2BX1 $T=1567220 1465750 0 0 $X=1567218 $Y=1465498
X87 339 15284 25 24 15260 NOR2BX1 $T=1569980 1421470 1 180 $X=1568140 $Y=1421218
X88 537 15280 25 24 15245 NOR2BX1 $T=1572740 1458370 0 180 $X=1570900 $Y=1454430
X89 383 15284 25 24 15332 NOR2BX1 $T=1571360 1421470 1 0 $X=1571358 $Y=1417530
X90 339 15335 25 24 15247 NOR2BX1 $T=1573200 1399330 0 180 $X=1571360 $Y=1395390
X91 537 15327 25 24 15194 NOR2BX1 $T=1573200 1487890 0 180 $X=1571360 $Y=1483950
X92 360 15323 25 24 15235 NOR2BX1 $T=1572740 1391950 1 0 $X=1572738 $Y=1388010
X93 339 15266 25 24 15322 NOR2BX1 $T=1572740 1465750 0 0 $X=1572738 $Y=1465498
X94 339 15323 25 24 15241 NOR2BX1 $T=1573200 1384570 1 0 $X=1573198 $Y=1380630
X95 391 15327 25 24 15337 NOR2BX1 $T=1573200 1473130 0 0 $X=1573198 $Y=1472878
X96 537 15132 25 24 15281 NOR2BX1 $T=1575040 1443610 0 180 $X=1573200 $Y=1439670
X97 10608 10669 25 24 16091 NOR2BX1 $T=1702460 1436230 0 0 $X=1702458 $Y=1435978
X98 10669 10608 25 24 16194 NOR2BX1 $T=1713040 1436230 1 0 $X=1713038 $Y=1432290
X99 9678 24 39 25 CLKBUFX3 $T=1091580 1443610 0 0 $X=1091578 $Y=1443358
X100 9902 24 9907 25 CLKBUFX3 $T=1103540 1450990 1 0 $X=1103538 $Y=1447050
X101 9994 24 10005 25 CLKBUFX3 $T=1112280 1443610 0 0 $X=1112278 $Y=1443358
X102 9920 24 102 25 CLKBUFX3 $T=1142640 1384570 0 0 $X=1142638 $Y=1384318
X103 10595 24 125 25 CLKBUFX3 $T=1161500 1362430 1 0 $X=1161498 $Y=1358490
X104 104 24 10126 25 CLKBUFX3 $T=1163340 1391950 0 0 $X=1163338 $Y=1391698
X105 10628 24 131 25 CLKBUFX3 $T=1166100 1369810 0 180 $X=1164260 $Y=1365870
X106 10582 24 135 25 CLKBUFX3 $T=1165640 1362430 1 0 $X=1165638 $Y=1358490
X107 10522 24 136 25 CLKBUFX3 $T=1166100 1355050 0 0 $X=1166098 $Y=1354798
X108 10645 24 137 25 CLKBUFX3 $T=1169320 1362430 1 0 $X=1169318 $Y=1358490
X109 10636 24 84 25 CLKBUFX3 $T=1172540 1487890 1 0 $X=1172538 $Y=1483950
X110 149 24 10803 25 CLKBUFX3 $T=1178060 1480510 1 0 $X=1178058 $Y=1476570
X111 10803 24 10810 25 CLKBUFX3 $T=1178060 1487890 1 0 $X=1178058 $Y=1483950
X112 10803 24 10469 25 CLKBUFX3 $T=1179900 1480510 1 180 $X=1178060 $Y=1480258
X113 10816 24 153 25 CLKBUFX3 $T=1179900 1362430 1 0 $X=1179898 $Y=1358490
X114 10803 24 10512 25 CLKBUFX3 $T=1182200 1487890 1 0 $X=1182198 $Y=1483950
X115 10512 24 10915 25 CLKBUFX3 $T=1182200 1524790 0 0 $X=1182198 $Y=1524538
X116 10512 24 11300 25 CLKBUFX3 $T=1208880 1532170 0 0 $X=1208878 $Y=1531918
X117 11305 24 200 25 CLKBUFX3 $T=1218080 1384570 1 0 $X=1218078 $Y=1380630
X118 11170 24 203 25 CLKBUFX3 $T=1219920 1384570 0 0 $X=1219918 $Y=1384318
X119 11487 24 10569 25 CLKBUFX3 $T=1231420 1532170 0 180 $X=1229580 $Y=1528230
X120 10279 24 164 25 CLKBUFX3 $T=1232340 1443610 0 0 $X=1232338 $Y=1443358
X121 10756 24 11692 25 CLKBUFX3 $T=1240160 1480510 1 0 $X=1240158 $Y=1476570
X122 11310 24 11794 25 CLKBUFX3 $T=1243380 1428850 1 0 $X=1243378 $Y=1424910
X123 10864 24 11804 25 CLKBUFX3 $T=1243840 1480510 1 0 $X=1243838 $Y=1476570
X124 11927 24 11907 25 CLKBUFX3 $T=1255800 1428850 1 180 $X=1253960 $Y=1428598
X125 11487 24 12054 25 CLKBUFX3 $T=1259940 1473130 1 0 $X=1259938 $Y=1469190
X126 12026 24 11869 25 CLKBUFX3 $T=1262240 1428850 0 180 $X=1260400 $Y=1424910
X127 12187 24 12071 25 CLKBUFX3 $T=1273280 1436230 0 180 $X=1271440 $Y=1432290
X128 10880 24 12253 25 CLKBUFX3 $T=1278340 1480510 1 0 $X=1278338 $Y=1476570
X129 12182 24 12224 25 CLKBUFX3 $T=1286160 1436230 0 180 $X=1284320 $Y=1432290
X130 12239 24 266 25 CLKBUFX3 $T=1289840 1399330 1 0 $X=1289838 $Y=1395390
X131 12364 24 12347 25 CLKBUFX3 $T=1290300 1377190 0 0 $X=1290298 $Y=1376938
X132 268 24 296 25 CLKBUFX3 $T=1293520 1399330 0 0 $X=1293518 $Y=1399078
X133 285 24 283 25 CLKBUFX3 $T=1293980 1458370 1 0 $X=1293978 $Y=1454430
X134 316 24 10062 25 CLKBUFX3 $T=1302720 1399330 0 180 $X=1300880 $Y=1395390
X135 276 24 294 25 CLKBUFX3 $T=1302260 1355050 1 0 $X=1302258 $Y=1351110
X136 316 24 268 25 CLKBUFX3 $T=1304100 1399330 0 0 $X=1304098 $Y=1399078
X137 316 24 288 25 CLKBUFX3 $T=1308700 1399330 1 0 $X=1308698 $Y=1395390
X138 329 24 12528 25 CLKBUFX3 $T=1312380 1355050 1 0 $X=1312378 $Y=1351110
X139 268 24 322 25 CLKBUFX3 $T=1312380 1399330 1 0 $X=1312378 $Y=1395390
X140 268 24 327 25 CLKBUFX3 $T=1312840 1391950 1 0 $X=1312838 $Y=1388010
X141 316 24 12404 25 CLKBUFX3 $T=1314220 1399330 0 0 $X=1314218 $Y=1399078
X142 12628 24 12330 25 CLKBUFX3 $T=1314680 1450990 0 0 $X=1314678 $Y=1450738
X143 268 24 321 25 CLKBUFX3 $T=1316520 1391950 1 0 $X=1316518 $Y=1388010
X144 333 24 12489 25 CLKBUFX3 $T=1316980 1369810 1 0 $X=1316978 $Y=1365870
X145 316 24 12641 25 CLKBUFX3 $T=1317900 1384570 1 0 $X=1317898 $Y=1380630
X146 12709 24 337 25 CLKBUFX3 $T=1322500 1399330 1 0 $X=1322498 $Y=1395390
X147 341 24 12525 25 CLKBUFX3 $T=1325260 1369810 0 180 $X=1323420 $Y=1365870
X148 316 24 348 25 CLKBUFX3 $T=1324340 1399330 1 0 $X=1324338 $Y=1395390
X149 39 24 347 25 CLKBUFX3 $T=1328940 1399330 0 0 $X=1328938 $Y=1399078
X150 355 24 12874 25 CLKBUFX3 $T=1330320 1355050 0 0 $X=1330318 $Y=1354798
X151 39 24 357 25 CLKBUFX3 $T=1331700 1399330 0 0 $X=1331698 $Y=1399078
X152 368 24 12726 25 CLKBUFX3 $T=1334460 1377190 0 0 $X=1334458 $Y=1376938
X153 39 24 358 25 CLKBUFX3 $T=1334920 1369810 0 0 $X=1334918 $Y=1369558
X154 39 24 374 25 CLKBUFX3 $T=1337220 1421470 1 0 $X=1337218 $Y=1417530
X155 39 24 360 25 CLKBUFX3 $T=1339060 1421470 0 0 $X=1339058 $Y=1421218
X156 39 24 382 25 CLKBUFX3 $T=1345500 1406710 1 0 $X=1345498 $Y=1402770
X157 39 24 383 25 CLKBUFX3 $T=1345500 1421470 1 0 $X=1345498 $Y=1417530
X158 369 24 12675 25 CLKBUFX3 $T=1346420 1355050 1 0 $X=1346418 $Y=1351110
X159 371 24 12806 25 CLKBUFX3 $T=1353780 1362430 1 0 $X=1353778 $Y=1358490
X160 39 24 386 25 CLKBUFX3 $T=1353780 1428850 0 0 $X=1353778 $Y=1428598
X161 12709 24 375 25 CLKBUFX3 $T=1358840 1399330 0 0 $X=1358838 $Y=1399078
X162 39 24 401 25 CLKBUFX3 $T=1362980 1428850 0 0 $X=1362978 $Y=1428598
X163 12559 24 403 25 CLKBUFX3 $T=1363440 1391950 0 0 $X=1363438 $Y=1391698
X164 12559 24 405 25 CLKBUFX3 $T=1365740 1384570 1 0 $X=1365738 $Y=1380630
X165 411 24 13241 25 CLKBUFX3 $T=1369420 1362430 1 0 $X=1369418 $Y=1358490
X166 316 24 13225 25 CLKBUFX3 $T=1369880 1384570 0 0 $X=1369878 $Y=1384318
X167 13298 24 12957 25 CLKBUFX3 $T=1371260 1561690 1 0 $X=1371258 $Y=1557750
X168 423 24 13312 25 CLKBUFX3 $T=1371720 1355050 0 0 $X=1371718 $Y=1354798
X169 12709 24 402 25 CLKBUFX3 $T=1373560 1399330 1 0 $X=1373558 $Y=1395390
X170 43 24 418 25 CLKBUFX3 $T=1379080 1391950 1 0 $X=1379078 $Y=1388010
X171 439 24 13313 25 CLKBUFX3 $T=1385520 1369810 0 0 $X=1385518 $Y=1369558
X172 316 24 431 25 CLKBUFX3 $T=1389200 1377190 0 0 $X=1389198 $Y=1376938
X173 438 24 13434 25 CLKBUFX3 $T=1397940 1362430 0 0 $X=1397938 $Y=1362178
X174 12709 24 381 25 CLKBUFX3 $T=1403000 1391950 1 180 $X=1401160 $Y=1391698
X175 316 24 455 25 CLKBUFX3 $T=1403000 1384570 1 0 $X=1402998 $Y=1380630
X176 12709 24 407 25 CLKBUFX3 $T=1403000 1414090 1 0 $X=1402998 $Y=1410150
X177 403 24 13143 25 CLKBUFX3 $T=1415420 1443610 1 0 $X=1415418 $Y=1439670
X178 463 24 13517 25 CLKBUFX3 $T=1419560 1369810 1 180 $X=1417720 $Y=1369558
X179 43 24 393 25 CLKBUFX3 $T=1419560 1450990 1 0 $X=1419558 $Y=1447050
X180 12709 24 469 25 CLKBUFX3 $T=1420020 1399330 0 0 $X=1420018 $Y=1399078
X181 295 24 472 25 CLKBUFX3 $T=1420940 1369810 1 0 $X=1420938 $Y=1365870
X182 274 24 13836 25 CLKBUFX3 $T=1421400 1450990 1 0 $X=1421398 $Y=1447050
X183 316 24 13723 25 CLKBUFX3 $T=1422320 1362430 0 0 $X=1422318 $Y=1362178
X184 299 24 13844 25 CLKBUFX3 $T=1423240 1406710 0 0 $X=1423238 $Y=1406458
X185 309 24 13850 25 CLKBUFX3 $T=1423700 1384570 1 0 $X=1423698 $Y=1380630
X186 12709 24 447 25 CLKBUFX3 $T=1423700 1399330 1 0 $X=1423698 $Y=1395390
X187 127 24 334 25 CLKBUFX3 $T=1423700 1436230 1 0 $X=1423698 $Y=1432290
X188 305 24 13877 25 CLKBUFX3 $T=1423700 1465750 0 0 $X=1423698 $Y=1465498
X189 127 24 12810 25 CLKBUFX3 $T=1423700 1480510 0 0 $X=1423698 $Y=1480258
X190 127 24 351 25 CLKBUFX3 $T=1425080 1473130 1 0 $X=1425078 $Y=1469190
X191 280 24 471 25 CLKBUFX3 $T=1427840 1355050 1 0 $X=1427838 $Y=1351110
X192 12709 24 477 25 CLKBUFX3 $T=1427840 1369810 0 0 $X=1427838 $Y=1369558
X193 43 24 410 25 CLKBUFX3 $T=1428760 1428850 0 0 $X=1428758 $Y=1428598
X194 298 24 13894 25 CLKBUFX3 $T=1428760 1502650 1 0 $X=1428758 $Y=1498710
X195 483 24 13885 25 CLKBUFX3 $T=1432440 1384570 1 0 $X=1432438 $Y=1380630
X196 311 24 13891 25 CLKBUFX3 $T=1432440 1399330 1 0 $X=1432438 $Y=1395390
X197 127 24 12724 25 CLKBUFX3 $T=1432440 1436230 1 0 $X=1432438 $Y=1432290
X198 12828 24 398 25 CLKBUFX3 $T=1432440 1443610 1 0 $X=1432438 $Y=1439670
X199 127 24 12718 25 CLKBUFX3 $T=1432440 1465750 0 0 $X=1432438 $Y=1465498
X200 476 24 486 25 CLKBUFX3 $T=1433360 1355050 1 0 $X=1433358 $Y=1351110
X201 127 24 12729 25 CLKBUFX3 $T=1433820 1428850 0 0 $X=1433818 $Y=1428598
X202 484 24 12735 25 CLKBUFX3 $T=1433820 1502650 1 0 $X=1433818 $Y=1498710
X203 43 24 396 25 CLKBUFX3 $T=1434280 1377190 0 0 $X=1434278 $Y=1376938
X204 12709 24 478 25 CLKBUFX3 $T=1434740 1406710 1 0 $X=1434738 $Y=1402770
X205 12709 24 475 25 CLKBUFX3 $T=1436580 1414090 0 0 $X=1436578 $Y=1413838
X206 488 24 13980 25 CLKBUFX3 $T=1440720 1391950 1 0 $X=1440718 $Y=1388010
X207 12709 24 480 25 CLKBUFX3 $T=1440720 1391950 0 0 $X=1440718 $Y=1391698
X208 284 24 14032 25 CLKBUFX3 $T=1440720 1539550 0 0 $X=1440718 $Y=1539298
X209 12709 24 494 25 CLKBUFX3 $T=1445780 1377190 1 0 $X=1445778 $Y=1373250
X210 12709 24 479 25 CLKBUFX3 $T=1449460 1391950 1 0 $X=1449458 $Y=1388010
X211 484 24 12788 25 CLKBUFX3 $T=1450380 1465750 0 0 $X=1450378 $Y=1465498
X212 484 24 12820 25 CLKBUFX3 $T=1451760 1436230 0 0 $X=1451758 $Y=1435978
X213 13294 24 13928 25 CLKBUFX3 $T=1455440 1436230 0 0 $X=1455438 $Y=1435978
X214 107 24 433 25 CLKBUFX3 $T=1456820 1406710 1 0 $X=1456818 $Y=1402770
X215 12709 24 496 25 CLKBUFX3 $T=1458200 1406710 0 0 $X=1458198 $Y=1406458
X216 308 24 14230 25 CLKBUFX3 $T=1459580 1532170 0 0 $X=1459578 $Y=1531918
X217 12709 24 491 25 CLKBUFX3 $T=1460960 1406710 1 0 $X=1460958 $Y=1402770
X218 313 24 14255 25 CLKBUFX3 $T=1461880 1517410 1 0 $X=1461878 $Y=1513470
X219 12709 24 493 25 CLKBUFX3 $T=1463260 1414090 1 0 $X=1463258 $Y=1410150
X220 12709 24 495 25 CLKBUFX3 $T=1465100 1391950 0 0 $X=1465098 $Y=1391698
X221 12709 24 502 25 CLKBUFX3 $T=1465100 1406710 1 0 $X=1465098 $Y=1402770
X222 12709 24 482 25 CLKBUFX3 $T=1466940 1406710 0 0 $X=1466938 $Y=1406458
X223 489 24 13932 25 CLKBUFX3 $T=1467400 1377190 1 0 $X=1467398 $Y=1373250
X224 127 24 512 25 CLKBUFX3 $T=1467860 1406710 1 0 $X=1467858 $Y=1402770
X225 12709 24 487 25 CLKBUFX3 $T=1468320 1414090 1 0 $X=1468318 $Y=1410150
X226 484 24 12733 25 CLKBUFX3 $T=1468320 1495270 0 0 $X=1468318 $Y=1495018
X227 316 24 457 25 CLKBUFX3 $T=1468780 1391950 0 0 $X=1468778 $Y=1391698
X228 512 24 12734 25 CLKBUFX3 $T=1471540 1465750 0 180 $X=1469700 $Y=1461810
X229 433 24 13107 25 CLKBUFX3 $T=1470160 1465750 0 0 $X=1470158 $Y=1465498
X230 505 24 13959 25 CLKBUFX3 $T=1475220 1391950 1 0 $X=1475218 $Y=1388010
X231 310 24 14356 25 CLKBUFX3 $T=1475220 1399330 1 0 $X=1475218 $Y=1395390
X232 312 24 14421 25 CLKBUFX3 $T=1475220 1428850 0 0 $X=1475218 $Y=1428598
X233 484 24 12790 25 CLKBUFX3 $T=1485800 1414090 1 0 $X=1485798 $Y=1410150
X234 301 24 14467 25 CLKBUFX3 $T=1487180 1546930 1 0 $X=1487178 $Y=1542990
X235 501 24 14131 25 CLKBUFX3 $T=1488100 1377190 1 0 $X=1488098 $Y=1373250
X236 509 24 14358 25 CLKBUFX3 $T=1489480 1377190 0 0 $X=1489478 $Y=1376938
X237 510 24 13996 25 CLKBUFX3 $T=1489940 1377190 1 0 $X=1489938 $Y=1373250
X238 300 24 14450 25 CLKBUFX3 $T=1489940 1480510 1 0 $X=1489938 $Y=1476570
X239 523 24 14168 25 CLKBUFX3 $T=1490860 1384570 1 0 $X=1490858 $Y=1380630
X240 520 24 14318 25 CLKBUFX3 $T=1491780 1377190 0 0 $X=1491778 $Y=1376938
X241 537 24 492 25 CLKBUFX3 $T=1508800 1369810 0 180 $X=1506960 $Y=1365870
X242 517 24 14273 25 CLKBUFX3 $T=1509260 1369810 1 0 $X=1509258 $Y=1365870
X243 537 24 485 25 CLKBUFX3 $T=1511560 1480510 1 180 $X=1509720 $Y=1480258
X244 288 24 504 25 CLKBUFX3 $T=1514780 1355050 0 0 $X=1514778 $Y=1354798
X245 84 24 537 25 CLKBUFX3 $T=1518920 1362430 1 0 $X=1518918 $Y=1358490
X246 13590 24 13948 25 CLKBUFX3 $T=1519380 1539550 1 0 $X=1519378 $Y=1535610
X247 288 24 519 25 CLKBUFX3 $T=1519840 1355050 0 0 $X=1519838 $Y=1354798
X248 288 24 539 25 CLKBUFX3 $T=1527200 1377190 0 0 $X=1527198 $Y=1376938
X249 288 24 521 25 CLKBUFX3 $T=1528120 1362430 1 0 $X=1528118 $Y=1358490
X250 484 24 345 25 CLKBUFX3 $T=1539160 1450990 0 180 $X=1537320 $Y=1447050
X251 529 24 14859 25 CLKBUFX3 $T=1537780 1362430 1 0 $X=1537778 $Y=1358490
X252 14659 24 14770 25 CLKBUFX3 $T=1541920 1391950 1 180 $X=1540080 $Y=1391698
X253 512 24 549 25 CLKBUFX3 $T=1543300 1369810 0 0 $X=1543298 $Y=1369558
X254 568 24 13590 25 CLKBUFX3 $T=1551580 1546930 1 0 $X=1551578 $Y=1542990
X255 12518 24 589 25 CLKBUFX3 $T=1571360 1355050 1 0 $X=1571358 $Y=1351110
X256 15334 24 15320 25 CLKBUFX3 $T=1592520 1399330 0 180 $X=1590680 $Y=1395390
X257 565 24 605 25 CLKBUFX3 $T=1597120 1369810 1 0 $X=1597118 $Y=1365870
X258 627 24 140 25 CLKBUFX3 $T=1661060 1694530 1 180 $X=1659220 $Y=1694278
X259 9673 9807 9673 24 9814 25 9839 OAI2BB2XL $T=1092960 1406710 0 0 $X=1092958 $Y=1406458
X260 9673 10019 9673 24 10023 25 10022 OAI2BB2XL $T=1111360 1414090 1 0 $X=1111358 $Y=1410150
X261 10146 10187 10126 24 10049 25 10168 OAI2BB2XL $T=1130680 1428850 1 180 $X=1127920 $Y=1428598
X262 10355 35 35 24 10366 25 10393 OAI2BB2XL $T=1144020 1421470 1 0 $X=1144018 $Y=1417530
X263 10246 35 35 24 10395 25 10385 OAI2BB2XL $T=1146780 1406710 0 0 $X=1146778 $Y=1406458
X264 10367 35 35 24 10509 25 10453 OAI2BB2XL $T=1155980 1421470 0 0 $X=1155978 $Y=1421218
X265 10629 10881 10881 24 10892 25 10754 OAI2BB2XL $T=1180820 1487890 0 0 $X=1180818 $Y=1487638
X266 10951 10892 10959 24 10951 25 10962 OAI2BB2XL $T=1188180 1487890 1 0 $X=1188178 $Y=1483950
X267 11645 10954 11252 24 266 25 12225 OAI2BB2XL $T=1272360 1384570 0 0 $X=1272358 $Y=1384318
X268 11638 10954 11252 24 270 25 12220 OAI2BB2XL $T=1276040 1377190 0 0 $X=1276038 $Y=1376938
X269 596 595 594 24 15330 25 15255 OAI2BB2XL $T=1583320 1369810 0 180 $X=1580560 $Y=1365870
X270 600 594 587 24 15388 25 15331 OAI2BB2XL $T=1589760 1377190 0 180 $X=1587000 $Y=1373250
X271 601 595 587 24 593 25 15412 OAI2BB2XL $T=1590680 1355050 1 180 $X=1587920 $Y=1354798
X272 602 595 594 24 15336 25 15345 OAI2BB2XL $T=1592520 1369810 1 180 $X=1589760 $Y=1369558
X273 607 594 587 24 15473 25 15494 OAI2BB2XL $T=1600800 1377190 0 180 $X=1598040 $Y=1373250
X274 611 594 606 24 609 25 608 OAI2BB2XL $T=1603560 1355050 0 180 $X=1600800 $Y=1351110
X275 613 594 595 24 15465 25 15545 OAI2BB2XL $T=1607700 1362430 0 180 $X=1604940 $Y=1358490
X276 612 594 595 24 15546 25 15544 OAI2BB2XL $T=1607700 1369810 1 180 $X=1604940 $Y=1369558
X277 614 595 594 24 15399 25 15470 OAI2BB2XL $T=1610000 1362430 1 180 $X=1607240 $Y=1362178
X278 621 594 606 24 620 25 619 OAI2BB2XL $T=1618280 1355050 0 180 $X=1615520 $Y=1351110
X279 622 594 595 24 15598 25 15596 OAI2BB2XL $T=1622420 1369810 1 180 $X=1619660 $Y=1369558
X280 623 594 606 24 15595 25 15648 OAI2BB2XL $T=1624720 1362430 1 180 $X=1621960 $Y=1362178
X281 626 594 606 24 616 25 15602 OAI2BB2XL $T=1627020 1355050 1 180 $X=1624260 $Y=1354798
X282 9682 43 24 25 CLKBUFX4 $T=1099400 1421470 0 0 $X=1099398 $Y=1421218
X283 9823 44 24 25 CLKBUFX4 $T=1104920 1421470 0 0 $X=1104918 $Y=1421218
X284 10122 74 24 25 CLKBUFX4 $T=1150920 1495270 0 0 $X=1150918 $Y=1495018
X285 39 344 24 25 CLKBUFX4 $T=1329860 1399330 1 0 $X=1329858 $Y=1395390
X286 39 391 24 25 CLKBUFX4 $T=1351940 1436230 1 0 $X=1351938 $Y=1432290
X287 624 149 24 25 CLKBUFX4 $T=1625640 1753570 1 180 $X=1623340 $Y=1753318
X288 9748 9747 9743 32 9683 9675 25 24 9674 SDFFRXL $T=1087900 1428850 0 180 $X=1076860 $Y=1424910
X289 9748 9749 9675 9741 9683 9680 25 24 9678 SDFFRXL $T=1088820 1443610 1 180 $X=1077780 $Y=1443358
X290 9748 9753 9680 9741 9683 9686 25 24 9682 SDFFRXL $T=1090660 1443610 0 180 $X=1079620 $Y=1439670
X291 9748 9755 9759 9741 9683 9841 25 24 9902 SDFFRXL $T=1089280 1458370 1 0 $X=1089278 $Y=1454430
X292 9911 9909 9838 32 9901 9803 25 24 9762 SDFFRXL $T=1102620 1377190 1 180 $X=1091580 $Y=1376938
X293 9748 9806 9686 9741 9683 9837 25 24 9994 SDFFRXL $T=1092040 1443610 1 0 $X=1092038 $Y=1439670
X294 9748 9921 9918 9741 9683 9826 25 24 9818 SDFFRXL $T=1105840 1473130 1 180 $X=1094800 $Y=1472878
X295 9748 9923 9919 32 9683 9743 25 24 9823 SDFFRXL $T=1106300 1428850 0 180 $X=1095260 $Y=1424910
X296 9748 9825 9837 9741 9901 9832 25 24 9810 SDFFRXL $T=1096640 1436230 1 0 $X=1096638 $Y=1432290
X297 9748 9835 9841 9741 9683 9918 25 24 9945 SDFFRXL $T=1097100 1465750 0 0 $X=1097098 $Y=1465498
X298 9911 9944 57 32 9901 9838 25 24 9819 SDFFRXL $T=1109060 1369810 1 180 $X=1098020 $Y=1369558
X299 9748 9991 9949 9741 9683 9759 25 24 9904 SDFFRXL $T=1111360 1458370 0 180 $X=1100320 $Y=1454430
X300 9748 10058 10049 32 9901 9919 25 24 58 SDFFRXL $T=1117800 1428850 0 180 $X=1106760 $Y=1424910
X301 9748 9951 9832 9741 10062 10070 25 24 10073 SDFFRXL $T=1108600 1436230 0 0 $X=1108598 $Y=1435978
X302 9911 10072 10069 32 75 62 25 24 9953 SDFFRXL $T=1120560 1355050 1 180 $X=1109520 $Y=1354798
X303 9952 10010 9826 9741 9683 10116 25 24 10007 SDFFRXL $T=1110900 1473130 0 0 $X=1110898 $Y=1472878
X304 9911 10113 10028 32 9901 10002 25 24 9816 SDFFRXL $T=1121940 1384570 0 180 $X=1110900 $Y=1380630
X305 9952 10017 10016 9741 10066 10119 25 24 10133 SDFFRXL $T=1111820 1517410 1 0 $X=1111818 $Y=1513470
X306 9952 10118 10114 9741 10066 10016 25 24 10011 SDFFRXL $T=1122860 1502650 1 180 $X=1111820 $Y=1502398
X307 9952 10128 10116 9741 9683 10026 25 24 10006 SDFFRXL $T=1123780 1480510 0 180 $X=1112740 $Y=1476570
X308 9911 10130 9803 32 9901 10028 25 24 9738 SDFFRXL $T=1124240 1377190 1 180 $X=1113200 $Y=1376938
X309 9952 10027 10026 9741 10066 10063 25 24 10155 SDFFRXL $T=1114120 1480510 0 0 $X=1114118 $Y=1480258
X310 9911 10141 10002 32 9901 10046 25 24 9677 SDFFRXL $T=1125160 1384570 1 180 $X=1114120 $Y=1384318
X311 9748 10051 10059 9741 9901 10136 25 24 91 SDFFRXL $T=1114580 1443610 0 0 $X=1114578 $Y=1443358
X312 9748 10147 10136 9741 9901 9949 25 24 70 SDFFRXL $T=1125620 1450990 1 180 $X=1114580 $Y=1450738
X313 9952 10057 10063 9741 10066 10132 25 24 10034 SDFFRXL $T=1115040 1487890 1 0 $X=1115038 $Y=1483950
X314 9911 10150 10142 32 9901 10055 25 24 9836 SDFFRXL $T=1126080 1399330 1 180 $X=1115040 $Y=1399078
X315 10154 10151 10055 32 10062 10056 25 24 72 SDFFRXL $T=1126080 1421470 0 180 $X=1115040 $Y=1417530
X316 9748 10168 10056 32 10062 10049 25 24 79 SDFFRXL $T=1128840 1428850 0 180 $X=1117800 $Y=1424910
X317 9952 10075 10132 9741 10066 10114 25 24 9995 SDFFRXL $T=1121020 1495270 1 0 $X=1121018 $Y=1491330
X318 9911 10240 10171 32 9901 10142 25 24 9831 SDFFRXL $T=1134820 1406710 1 180 $X=1123780 $Y=1406458
X319 9911 10252 10046 32 9901 10165 25 24 9737 SDFFRXL $T=1137120 1384570 1 180 $X=1126080 $Y=1384318
X320 9911 10167 10165 32 9901 10253 25 24 10025 SDFFRXL $T=1126540 1391950 0 0 $X=1126538 $Y=1391698
X321 9911 10257 10253 32 9901 10170 25 24 9899 SDFFRXL $T=1138040 1399330 0 180 $X=1127000 $Y=1395390
X322 9911 10258 10170 32 9901 10171 25 24 9829 SDFFRXL $T=1138040 1406710 0 180 $X=1127000 $Y=1402770
X323 9748 10259 10236 9741 9901 10059 25 24 10135 SDFFRXL $T=1138040 1450990 1 180 $X=1127000 $Y=1450738
X324 9952 10175 10119 9741 10066 10228 25 24 10291 SDFFRXL $T=1127460 1517410 1 0 $X=1127458 $Y=1513470
X325 9952 10189 10228 9741 10066 10278 25 24 10283 SDFFRXL $T=1129300 1510030 1 0 $X=1129298 $Y=1506090
X326 10154 10276 10269 32 10062 10222 25 24 93 SDFFRXL $T=1140800 1428850 0 180 $X=1129760 $Y=1424910
X327 9748 10229 10070 9741 10062 10269 25 24 97 SDFFRXL $T=1130680 1436230 0 0 $X=1130678 $Y=1435978
X328 9911 10296 10239 32 10062 10233 25 24 9813 SDFFRXL $T=1142180 1377190 1 180 $X=1131140 $Y=1376938
X329 9748 10235 10222 32 10062 10342 25 24 10355 SDFFRXL $T=1131600 1421470 1 0 $X=1131598 $Y=1417530
X330 9748 10337 10288 9741 9901 10236 25 24 10223 SDFFRXL $T=1142640 1450990 0 180 $X=1131600 $Y=1447050
X331 9911 10286 10250 32 10062 10239 25 24 9842 SDFFRXL $T=1143560 1391950 0 180 $X=1132520 $Y=1388010
X332 10154 10357 10342 32 9901 10250 25 24 10246 SDFFRXL $T=1145860 1406710 1 180 $X=1134820 $Y=1406458
X333 9952 10347 10278 9741 10066 10381 25 24 10470 SDFFRXL $T=1141260 1510030 1 0 $X=1141258 $Y=1506090
X334 9911 10479 10233 32 10062 10363 25 24 9808 SDFFRXL $T=1155060 1369810 1 180 $X=1144020 $Y=1369558
X335 10241 10480 10399 9741 9901 10358 25 24 106 SDFFRXL $T=1155060 1443610 0 180 $X=1144020 $Y=1439670
X336 9952 10368 10381 9741 10066 10482 25 24 10491 SDFFRXL $T=1144940 1502650 0 0 $X=1144938 $Y=1502398
X337 10154 10385 10392 32 112 10395 25 24 10507 SDFFRXL $T=1146320 1406710 1 0 $X=1146318 $Y=1402770
X338 10241 10379 10401 9741 10062 10361 25 24 10510 SDFFRXL $T=1147240 1428850 0 0 $X=1147238 $Y=1428598
X339 10241 10500 10358 9741 9901 10288 25 24 10388 SDFFRXL $T=1158280 1443610 1 180 $X=1147240 $Y=1443358
X340 9911 10360 10398 32 116 10372 25 24 123 SDFFRXL $T=1148620 1384570 0 0 $X=1148618 $Y=1384318
X341 9911 10445 10372 32 116 10484 25 24 126 SDFFRXL $T=1148620 1391950 1 0 $X=1148618 $Y=1388010
X342 10154 10393 115 32 112 10366 25 24 10593 SDFFRXL $T=1148620 1421470 1 0 $X=1148618 $Y=1417530
X343 9952 10448 10458 9741 10066 10521 25 24 10581 SDFFRXL $T=1148620 1517410 1 0 $X=1148618 $Y=1513470
X344 10241 10394 10509 32 10062 10401 25 24 10367 SDFFRXL $T=1159660 1428850 0 180 $X=1148620 $Y=1424910
X345 10241 10519 10510 9741 10062 10446 25 24 10399 SDFFRXL $T=1159660 1436230 1 180 $X=1148620 $Y=1435978
X346 10154 10452 10462 32 10469 10518 25 24 10589 SDFFRXL $T=1149080 1414090 1 0 $X=1149078 $Y=1410150
X347 10154 10453 10395 32 112 10509 25 24 10577 SDFFRXL $T=1149080 1414090 0 0 $X=1149078 $Y=1413838
X348 9911 10384 10397 32 116 10398 25 24 130 SDFFRXL $T=1149540 1384570 1 0 $X=1149538 $Y=1380630
X349 9911 10383 10517 32 116 10397 25 24 113 SDFFRXL $T=1160580 1377190 0 180 $X=1149540 $Y=1373250
X350 10154 10533 10484 32 116 10392 25 24 114 SDFFRXL $T=1160580 1399330 0 180 $X=1149540 $Y=1395390
X351 10569 10536 10521 9741 10512 10459 25 24 9998 SDFFRXL $T=1160580 1524790 1 180 $X=1149540 $Y=1524538
X352 9911 10464 10363 32 116 10517 25 24 129 SDFFRXL $T=1150460 1369810 1 0 $X=1150458 $Y=1365870
X353 9952 10476 10482 9741 10066 10458 25 24 10600 SDFFRXL $T=1152300 1510030 1 0 $X=1152298 $Y=1506090
X354 10154 10508 10518 32 10469 10642 25 24 10648 SDFFRXL $T=1156440 1406710 0 0 $X=1156438 $Y=1406458
X355 10241 10535 10534 9741 116 10664 25 24 10645 SDFFRXL $T=1158280 1450990 1 0 $X=1158278 $Y=1447050
X356 10241 10657 10590 9741 116 10534 25 24 10522 SDFFRXL $T=1169320 1443610 1 180 $X=1158280 $Y=1443358
X357 10241 10677 10670 9741 116 10590 25 24 10582 SDFFRXL $T=1171620 1458370 1 180 $X=1160580 $Y=1458118
X358 10154 10713 10598 10663 10469 10462 25 24 10588 SDFFRXL $T=1172080 1414090 1 180 $X=1161040 $Y=1413838
X359 10241 10717 10643 10663 10469 10598 25 24 10591 SDFFRXL $T=1172540 1428850 0 180 $X=1161500 $Y=1424910
X360 10569 10729 10651 9741 10066 10609 25 24 10511 SDFFRXL $T=1173920 1517410 1 180 $X=1162880 $Y=1517158
X361 10569 10611 10625 9741 9683 10670 25 24 10636 SDFFRXL $T=1163340 1487890 0 0 $X=1163338 $Y=1487638
X362 9952 10633 10609 9741 10066 10744 25 24 10763 SDFFRXL $T=1164720 1517410 1 0 $X=1164718 $Y=1513470
X363 10569 10634 10459 9741 10512 10745 25 24 10122 SDFFRXL $T=1164720 1524790 0 0 $X=1164718 $Y=1524538
X364 10569 10754 10738 9741 10512 10625 25 24 10629 SDFFRXL $T=1176220 1495270 0 180 $X=1165180 $Y=1491330
X365 10569 10626 10649 9741 10512 10738 25 24 10596 SDFFRXL $T=1165640 1495270 0 0 $X=1165638 $Y=1495018
X366 10241 10761 10710 9741 10469 10643 25 24 10635 SDFFRXL $T=1176680 1436230 0 180 $X=1165640 $Y=1432290
X367 10569 10769 10650 9741 10066 10649 25 24 10614 SDFFRXL $T=1177140 1502650 1 180 $X=1166100 $Y=1502398
X368 10569 10770 10744 9741 10066 10650 25 24 10505 SDFFRXL $T=1177140 1510030 0 180 $X=1166100 $Y=1506090
X369 10569 10771 10755 9741 10066 10651 25 24 10583 SDFFRXL $T=1177140 1524790 0 180 $X=1166100 $Y=1520850
X370 10241 10711 10664 9741 116 10808 25 24 10816 SDFFRXL $T=1169320 1450990 1 0 $X=1169318 $Y=1447050
X371 10241 10807 10799 9741 10469 10710 25 24 10671 SDFFRXL $T=1180360 1443610 1 180 $X=1169320 $Y=1443358
X372 10241 10950 10900 9741 10469 10799 25 24 10802 SDFFRXL $T=1189560 1465750 0 180 $X=1178520 $Y=1461810
X373 10569 10851 10745 9741 10512 10755 25 24 10929 SDFFRXL $T=1179440 1532170 1 0 $X=1179438 $Y=1528230
X374 11028 11029 10918 9741 10469 10900 25 24 10894 SDFFRXL $T=1193700 1473130 1 180 $X=1182660 $Y=1472878
X375 10154 11020 161 10663 10810 10902 25 24 10742 SDFFRXL $T=1194160 1391950 0 180 $X=1183120 $Y=1388010
X376 11028 10898 160 10663 10810 10914 25 24 10798 SDFFRXL $T=1194620 1399330 0 180 $X=1183580 $Y=1395390
X377 10154 10855 10928 10663 10915 11017 25 24 10762 SDFFRXL $T=1184040 1414090 0 0 $X=1184038 $Y=1413838
X378 10154 10944 10642 10663 10469 11066 25 24 11082 SDFFRXL $T=1186800 1414090 1 0 $X=1186798 $Y=1410150
X379 11028 11072 11066 10663 10469 10928 25 24 10938 SDFFRXL $T=1198300 1421470 0 180 $X=1187260 $Y=1417530
X380 11028 11033 168 10663 10810 11170 25 24 11178 SDFFRXL $T=1191860 1391950 0 0 $X=1191858 $Y=1391698
X381 11028 11195 11185 10663 10512 11067 25 24 11060 SDFFRXL $T=1206120 1495270 1 180 $X=1195080 $Y=1495018
X382 10241 11061 11083 10663 10915 11206 25 24 10737 SDFFRXL $T=1196000 1421470 0 0 $X=1195998 $Y=1421218
X383 10569 11076 11092 10663 10512 11185 25 24 11235 SDFFRXL $T=1196460 1502650 0 0 $X=1196458 $Y=1502398
X384 10569 11198 11214 10663 10512 11092 25 24 11071 SDFFRXL $T=1208880 1532170 1 180 $X=1197840 $Y=1531918
X385 11028 11167 11067 10663 10469 11204 25 24 11260 SDFFRXL $T=1200140 1487890 1 0 $X=1200138 $Y=1483950
X386 10241 11250 11234 10663 10469 11083 25 24 11126 SDFFRXL $T=1211180 1421470 0 180 $X=1200140 $Y=1417530
X387 10241 11099 187 10663 10915 11166 25 24 10887 SDFFRXL $T=1211180 1443610 0 180 $X=1200140 $Y=1439670
X388 11028 11183 180 10663 10810 11305 25 24 11313 SDFFRXL $T=1202900 1391950 0 0 $X=1202898 $Y=1391698
X389 11028 11379 201 10663 10915 11310 25 24 11203 SDFFRXL $T=1224060 1443610 0 180 $X=1213020 $Y=1439670
X390 10241 11443 202 10663 10915 11311 25 24 11227 SDFFRXL $T=1224060 1458370 1 180 $X=1213020 $Y=1458118
X391 11028 11449 11437 10663 11300 11234 25 24 11314 SDFFRXL $T=1224520 1421470 0 180 $X=1213480 $Y=1417530
X392 10569 11481 11470 10663 10915 11356 25 24 11317 SDFFRXL $T=1226820 1517410 1 180 $X=1215780 $Y=1517158
X393 11487 11476 11471 10663 11300 11214 25 24 11346 SDFFRXL $T=1226820 1532170 1 180 $X=1215780 $Y=1531918
X394 11028 11538 208 10663 10915 11438 25 24 11362 SDFFRXL $T=1232340 1480510 1 180 $X=1221300 $Y=1480258
X395 11028 11461 211 10663 10915 11480 25 24 11316 SDFFRXL $T=1235560 1502650 0 180 $X=1224520 $Y=1498710
X396 11487 11532 11542 10663 11300 11471 25 24 11772 SDFFRXL $T=1229580 1539550 0 0 $X=1229578 $Y=1539298
X397 11487 11658 11674 10663 11300 11542 25 24 11539 SDFFRXL $T=1242000 1539550 0 180 $X=1230960 $Y=1535610
X398 11028 11501 210 10663 10810 11687 25 24 11647 SDFFRXL $T=1231420 1399330 1 0 $X=1231418 $Y=1395390
X399 11487 11640 217 10663 10915 11777 25 24 11690 SDFFRXL $T=1235100 1495270 1 0 $X=1235098 $Y=1491330
X400 11028 11668 11755 10663 11300 11437 25 24 11624 SDFFRXL $T=1246140 1421470 1 180 $X=1235100 $Y=1421218
X401 10154 11656 218 10663 11300 11792 25 24 11775 SDFFRXL $T=1236940 1384570 0 0 $X=1236938 $Y=1384318
X402 224 225 11789 229 230 11810 25 24 242 SDFFRXL $T=1244760 1369810 0 0 $X=1244758 $Y=1369558
X403 224 223 227 229 230 240 25 24 243 SDFFRXL $T=1245220 1355050 0 0 $X=1245218 $Y=1354798
X404 11487 11796 11806 10663 10915 11942 25 24 11918 SDFFRXL $T=1246600 1495270 0 0 $X=1246598 $Y=1495018
X405 224 11899 11912 229 230 11789 25 24 226 SDFFRXL $T=1257640 1369810 0 180 $X=1246600 $Y=1365870
X406 224 11773 11810 229 230 11914 25 24 237 SDFFRXL $T=1247060 1377190 1 0 $X=1247058 $Y=1373250
X407 11487 11893 11903 10663 11300 11674 25 24 11803 SDFFRXL $T=1259020 1539550 0 180 $X=1247980 $Y=1535610
X408 224 11868 233 229 11300 11917 25 24 11925 SDFFRXL $T=1248440 1391950 0 0 $X=1248438 $Y=1391698
X409 11874 11881 10808 10663 10915 11954 25 24 11920 SDFFRXL $T=1249360 1443610 0 0 $X=1249358 $Y=1443358
X410 11874 11927 11955 10663 10810 11755 25 24 11811 SDFFRXL $T=1260400 1443610 0 180 $X=1249360 $Y=1439670
X411 11487 11943 12013 11960 11300 11903 25 24 11895 SDFFRXL $T=1262240 1539550 1 180 $X=1251200 $Y=1539298
X412 11028 11905 11914 10663 11300 12025 25 24 12033 SDFFRXL $T=1251660 1414090 1 0 $X=1251658 $Y=1410150
X413 11487 11771 12017 11960 10915 11902 25 24 11739 SDFFRXL $T=1262700 1495270 0 180 $X=1251660 $Y=1491330
X414 11028 11913 11920 229 11300 12040 25 24 12117 SDFFRXL $T=1252580 1399330 1 0 $X=1252578 $Y=1395390
X415 11874 11915 11922 10663 10062 12034 25 24 12046 SDFFRXL $T=1252580 1450990 1 0 $X=1252578 $Y=1447050
X416 224 253 11945 229 230 11912 25 24 239 SDFFRXL $T=1264080 1362430 0 180 $X=1253040 $Y=1358490
X417 224 11924 11934 229 230 12052 25 24 254 SDFFRXL $T=1253960 1362430 0 0 $X=1253958 $Y=1362178
X418 224 11798 12045 229 230 11934 25 24 244 SDFFRXL $T=1266840 1369810 1 180 $X=1255800 $Y=1369558
X419 224 257 12052 229 230 11945 25 24 246 SDFFRXL $T=1267300 1355050 1 180 $X=1256260 $Y=1354798
X420 224 249 12171 229 230 12045 25 24 252 SDFFRXL $T=1273280 1377190 0 180 $X=1262240 $Y=1373250
X421 11874 12182 12064 12113 11300 11955 25 24 12036 SDFFRXL $T=1273280 1436230 1 180 $X=1262240 $Y=1435978
X422 11487 12103 12174 11960 11300 12013 25 24 12037 SDFFRXL $T=1273280 1539550 1 180 $X=1262240 $Y=1539298
X423 11028 12055 12025 229 11300 12175 25 24 12208 SDFFRXL $T=1264080 1414090 1 0 $X=1264078 $Y=1410150
X424 11487 12058 12066 11960 10915 12207 25 24 12173 SDFFRXL $T=1264080 1510030 1 0 $X=1264078 $Y=1506090
X425 224 267 265 229 258 256 25 24 255 SDFFRXL $T=1276040 1355050 0 180 $X=1265000 $Y=1351110
X426 11874 11873 12198 12113 11300 12064 25 24 12060 SDFFRXL $T=1276040 1428850 1 180 $X=1265000 $Y=1428598
X427 224 12112 12167 229 10810 12239 25 24 12230 SDFFRXL $T=1268680 1406710 1 0 $X=1268678 $Y=1402770
X428 224 11877 12226 229 230 12111 25 24 259 SDFFRXL $T=1279720 1362430 1 180 $X=1268680 $Y=1362178
X429 11874 12236 12227 12113 268 12114 25 24 12102 SDFFRXL $T=1279720 1450990 0 180 $X=1268680 $Y=1447050
X430 11487 12057 12232 12113 10915 12115 25 24 12014 SDFFRXL $T=1280180 1487890 1 180 $X=1269140 $Y=1487638
X431 11028 11957 12175 12113 11300 12188 25 24 12314 SDFFRXL $T=1269600 1421470 1 0 $X=1269598 $Y=1417530
X432 224 11675 12111 229 230 12249 25 24 273 SDFFRXL $T=1270060 1369810 1 0 $X=1270058 $Y=1365870
X433 11487 12099 245 11960 11300 12211 25 24 12322 SDFFRXL $T=1270060 1532170 1 0 $X=1270058 $Y=1528230
X434 11028 12116 264 229 11300 12313 25 24 12053 SDFFRXL $T=1270520 1391950 1 0 $X=1270518 $Y=1388010
X435 11874 12181 12188 12113 11300 12198 25 24 12327 SDFFRXL $T=1270980 1428850 1 0 $X=1270978 $Y=1424910
X436 224 11894 12249 229 230 12171 25 24 261 SDFFRXL $T=1282020 1369810 1 180 $X=1270980 $Y=1369558
X437 11487 12080 12211 11960 11300 12174 25 24 12343 SDFFRXL $T=1273280 1539550 0 0 $X=1273278 $Y=1539298
X438 11874 12333 12102 12113 10915 12205 25 24 12167 SDFFRXL $T=1284320 1436230 1 180 $X=1273280 $Y=1435978
X439 12054 12406 12403 12113 288 12317 25 24 12232 SDFFRXL $T=1291220 1480510 0 180 $X=1280180 $Y=1476570
X440 12411 12409 12379 11960 288 12318 25 24 12066 SDFFRXL $T=1291220 1517410 0 180 $X=1280180 $Y=1513470
X441 12054 12337 281 12113 288 12466 25 24 12339 SDFFRXL $T=1282480 1487890 1 0 $X=1282478 $Y=1483950
X442 11487 12340 286 11960 288 12472 25 24 12361 SDFFRXL $T=1282940 1502650 0 0 $X=1282938 $Y=1502398
X443 289 12407 12470 229 268 12355 25 24 12348 SDFFRXL $T=1295360 1369810 1 180 $X=1284320 $Y=1369558
X444 12478 12475 292 229 288 12356 25 24 12350 SDFFRXL $T=1295360 1414090 0 180 $X=1284320 $Y=1410150
X445 289 12376 12350 229 149 12412 25 24 12470 SDFFRXL $T=1285700 1391950 0 0 $X=1285698 $Y=1391698
X446 12411 12494 12483 11960 288 12386 25 24 12379 SDFFRXL $T=1297660 1510030 1 180 $X=1286620 $Y=1509778
X447 12054 12393 12361 11960 288 12504 25 24 12177 SDFFRXL $T=1287080 1495270 1 0 $X=1287078 $Y=1491330
X448 289 12394 293 229 288 306 25 24 12226 SDFFRXL $T=1287540 1362430 0 0 $X=1287538 $Y=1362178
X449 289 12396 12336 229 268 12509 25 24 12578 SDFFRXL $T=1287540 1377190 1 0 $X=1287538 $Y=1373250
X450 11874 12401 12369 12113 268 12481 25 24 12408 SDFFRXL $T=1288000 1428850 0 0 $X=1287998 $Y=1428598
X451 11874 12402 12408 12113 288 12510 25 24 12392 SDFFRXL $T=1288000 1436230 0 0 $X=1287998 $Y=1435978
X452 12054 12484 12339 12113 288 12465 25 24 12463 SDFFRXL $T=1302260 1480510 0 180 $X=1291220 $Y=1476570
X453 318 12580 317 229 149 10069 25 24 12476 SDFFRXL $T=1304560 1355050 1 180 $X=1293520 $Y=1354798
X454 12411 12624 12618 11960 288 12519 25 24 12483 SDFFRXL $T=1308700 1510030 1 180 $X=1297660 $Y=1509778
X455 565 15255 15234 586 75 15330 25 24 590 SDFFRXL $T=1564460 1369810 1 0 $X=1564458 $Y=1365870
X456 565 15331 15336 586 75 15388 25 24 597 SDFFRXL $T=1574120 1362430 1 0 $X=1574118 $Y=1358490
X457 565 15345 15330 586 75 15336 25 24 599 SDFFRXL $T=1577340 1369810 0 0 $X=1577338 $Y=1369558
X458 565 15412 15388 586 75 593 25 24 592 SDFFRXL $T=1591600 1355050 0 180 $X=1580560 $Y=1351110
X459 605 15470 15465 586 75 15399 25 24 598 SDFFRXL $T=1596200 1362430 0 180 $X=1585160 $Y=1358490
X460 605 15494 15399 586 75 15473 25 24 603 SDFFRXL $T=1605400 1362430 1 180 $X=1594360 $Y=1362178
X461 605 15545 609 586 610 15465 25 24 604 SDFFRXL $T=1610000 1355050 1 180 $X=1598960 $Y=1354798
X462 605 15544 15473 586 610 15546 25 24 617 SDFFRXL $T=1603100 1369810 1 0 $X=1603098 $Y=1365870
X463 605 15602 15595 586 610 616 25 24 615 SDFFRXL $T=1622880 1355050 1 180 $X=1611840 $Y=1354798
X464 605 15648 15598 586 610 15595 25 24 618 SDFFRXL $T=1626560 1362430 0 180 $X=1615520 $Y=1358490
X465 605 15596 15546 586 610 15598 25 24 625 SDFFRXL $T=1615980 1369810 1 0 $X=1615978 $Y=1365870
X466 9952 24 9748 25 CLKBUFX2 $T=1109060 1473130 0 0 $X=1109058 $Y=1472878
X467 10135 24 86 25 CLKBUFX2 $T=1124240 1384570 0 180 $X=1122400 $Y=1380630
X468 94 24 10033 25 CLKBUFX2 $T=1129300 1355050 1 0 $X=1129298 $Y=1351110
X469 9953 24 10137 25 CLKBUFX2 $T=1129300 1355050 0 0 $X=1129298 $Y=1354798
X470 9748 24 10241 25 CLKBUFX2 $T=1132060 1428850 0 0 $X=1132058 $Y=1428598
X471 10062 24 9901 25 CLKBUFX2 $T=1138960 1384570 0 0 $X=1138958 $Y=1384318
X472 10154 24 9911 25 CLKBUFX2 $T=1144480 1406710 1 0 $X=1144478 $Y=1402770
X473 10126 24 89 25 CLKBUFX2 $T=1148160 1391950 0 0 $X=1148158 $Y=1391698
X474 10577 24 10608 25 CLKBUFX2 $T=1161500 1436230 1 0 $X=1161498 $Y=1432290
X475 10578 24 9805 25 CLKBUFX2 $T=1162420 1502650 1 0 $X=1162418 $Y=1498710
X476 10593 24 10669 25 CLKBUFX2 $T=1162880 1428850 0 0 $X=1162878 $Y=1428598
X477 10387 24 9830 25 CLKBUFX2 $T=1164720 1502650 1 0 $X=1164718 $Y=1498710
X478 10661 24 138 25 CLKBUFX2 $T=1167940 1377190 1 0 $X=1167938 $Y=1373250
X479 10662 24 139 25 CLKBUFX2 $T=1170240 1355050 0 0 $X=1170238 $Y=1354798
X480 10716 24 147 25 CLKBUFX2 $T=1174380 1362430 0 0 $X=1174378 $Y=1362178
X481 10569 24 9952 25 CLKBUFX2 $T=1175760 1517410 1 0 $X=1175758 $Y=1513470
X482 10794 24 148 25 CLKBUFX2 $T=1178520 1384570 0 0 $X=1178518 $Y=1384318
X483 10721 24 152 25 CLKBUFX2 $T=1179440 1362430 0 0 $X=1179438 $Y=1362178
X484 10469 24 9683 25 CLKBUFX2 $T=1179900 1480510 0 0 $X=1179898 $Y=1480258
X485 10810 24 10066 25 CLKBUFX2 $T=1179900 1487890 1 0 $X=1179898 $Y=1483950
X486 10882 24 10371 25 CLKBUFX2 $T=1183120 1495270 1 180 $X=1181280 $Y=1495018
X487 10897 24 150 25 CLKBUFX2 $T=1182660 1384570 0 0 $X=1182658 $Y=1384318
X488 10902 24 154 25 CLKBUFX2 $T=1183120 1384570 1 0 $X=1183118 $Y=1380630
X489 10929 24 10460 25 CLKBUFX2 $T=1186800 1524790 1 180 $X=1184960 $Y=1524538
X490 11075 24 176 25 CLKBUFX2 $T=1196920 1391950 1 0 $X=1196918 $Y=1388010
X491 11079 24 179 25 CLKBUFX2 $T=1202900 1369810 1 0 $X=1202898 $Y=1365870
X492 10952 24 10760 25 CLKBUFX2 $T=1202900 1480510 1 0 $X=1202898 $Y=1476570
X493 11098 24 11249 25 CLKBUFX2 $T=1206580 1436230 0 0 $X=1206578 $Y=1435978
X494 11188 24 190 25 CLKBUFX2 $T=1207040 1362430 1 0 $X=1207038 $Y=1358490
X495 11163 24 191 25 CLKBUFX2 $T=1208420 1391950 1 0 $X=1208418 $Y=1388010
X496 10801 24 11321 25 CLKBUFX2 $T=1215780 1428850 0 0 $X=1215778 $Y=1428598
X497 11393 24 10925 25 CLKBUFX2 $T=1220380 1399330 0 0 $X=1220378 $Y=1399078
X498 11308 24 11486 25 CLKBUFX2 $T=1220840 1480510 1 0 $X=1220838 $Y=1476570
X499 11430 24 11496 25 CLKBUFX2 $T=1224520 1465750 1 0 $X=1224518 $Y=1461810
X500 11369 24 11530 25 CLKBUFX2 $T=1226360 1495270 1 0 $X=1226358 $Y=1491330
X501 11580 24 10954 25 CLKBUFX2 $T=1232800 1450990 1 0 $X=1232798 $Y=1447050
X502 11583 24 178 25 CLKBUFX2 $T=1233260 1362430 0 0 $X=1233258 $Y=1362178
X503 11105 24 10952 25 CLKBUFX2 $T=1236020 1480510 0 0 $X=1236018 $Y=1480258
X504 11179 24 162 25 CLKBUFX2 $T=1241540 1428850 1 0 $X=1241538 $Y=1424910
X505 224 24 10154 25 CLKBUFX2 $T=1247060 1391950 1 0 $X=1247058 $Y=1388010
X506 11736 24 231 25 CLKBUFX2 $T=1247980 1384570 1 0 $X=1247978 $Y=1380630
X507 11687 24 236 25 CLKBUFX2 $T=1249820 1399330 1 0 $X=1249818 $Y=1395390
X508 11917 24 11871 25 CLKBUFX2 $T=1254880 1391950 0 180 $X=1253040 $Y=1388010
X509 11920 24 11965 25 CLKBUFX2 $T=1254880 1428850 1 0 $X=1254878 $Y=1424910
X510 11327 24 10899 25 CLKBUFX2 $T=1256260 1436230 1 0 $X=1256258 $Y=1432290
X511 11942 24 12056 25 CLKBUFX2 $T=1259020 1487890 1 0 $X=1259018 $Y=1483950
X512 12016 24 248 25 CLKBUFX2 $T=1261320 1377190 0 180 $X=1259480 $Y=1373250
X513 11874 24 11028 25 CLKBUFX2 $T=1269140 1428850 1 0 $X=1269138 $Y=1424910
X514 11487 24 224 25 CLKBUFX2 $T=1269140 1473130 1 0 $X=1269138 $Y=1469190
X515 12167 24 12334 25 CLKBUFX2 $T=1276040 1443610 1 0 $X=1276038 $Y=1439670
X516 12054 24 11874 25 CLKBUFX2 $T=1289380 1473130 1 0 $X=1289378 $Y=1469190
X517 12476 24 12518 25 CLKBUFX2 $T=1293980 1362430 1 0 $X=1293978 $Y=1358490
X518 12347 24 314 25 CLKBUFX2 $T=1295820 1377190 0 0 $X=1295818 $Y=1376938
X519 12330 24 279 25 CLKBUFX2 $T=1297660 1414090 0 0 $X=1297658 $Y=1413838
X520 12253 24 275 25 CLKBUFX2 $T=1298580 1391950 1 0 $X=1298578 $Y=1388010
X521 12366 24 277 25 CLKBUFX2 $T=1303180 1391950 1 0 $X=1303178 $Y=1388010
X522 10062 24 324 25 CLKBUFX2 $T=1306400 1399330 1 0 $X=1306398 $Y=1395390
X523 12404 24 325 25 CLKBUFX2 $T=1309160 1399330 0 0 $X=1309158 $Y=1399078
X524 12411 24 12370 25 CLKBUFX2 $T=1312840 1517410 1 0 $X=1312838 $Y=1513470
X525 12528 24 330 25 CLKBUFX2 $T=1314220 1355050 1 0 $X=1314218 $Y=1351110
X526 268 24 12709 25 CLKBUFX2 $T=1314220 1399330 1 0 $X=1314218 $Y=1395390
X527 12489 24 336 25 CLKBUFX2 $T=1318820 1369810 1 0 $X=1318818 $Y=1365870
X528 12525 24 346 25 CLKBUFX2 $T=1325260 1369810 1 0 $X=1325258 $Y=1365870
X529 12874 24 363 25 CLKBUFX2 $T=1332160 1355050 0 0 $X=1332158 $Y=1354798
X530 12411 24 12597 25 CLKBUFX2 $T=1332620 1510030 0 0 $X=1332618 $Y=1509778
X531 365 24 12828 25 CLKBUFX2 $T=1333540 1399330 0 0 $X=1333538 $Y=1399078
X532 366 24 12478 25 CLKBUFX2 $T=1334000 1399330 1 0 $X=1333998 $Y=1395390
X533 12726 24 372 25 CLKBUFX2 $T=1336300 1377190 0 0 $X=1336298 $Y=1376938
X534 12957 24 12411 25 CLKBUFX2 $T=1339060 1554310 1 0 $X=1339058 $Y=1550370
X535 12641 24 380 25 CLKBUFX2 $T=1347340 1406710 1 0 $X=1347338 $Y=1402770
X536 12675 24 385 25 CLKBUFX2 $T=1348260 1355050 1 0 $X=1348258 $Y=1351110
X537 12806 24 390 25 CLKBUFX2 $T=1351940 1362430 1 0 $X=1351938 $Y=1358490
X538 13241 24 427 25 CLKBUFX2 $T=1371260 1362430 1 0 $X=1371258 $Y=1358490
X539 13312 24 434 25 CLKBUFX2 $T=1374480 1355050 0 0 $X=1374478 $Y=1354798
X540 13225 24 435 25 CLKBUFX2 $T=1377700 1369810 1 0 $X=1377698 $Y=1365870
X541 13272 24 12942 25 CLKBUFX2 $T=1385060 1428850 1 0 $X=1385058 $Y=1424910
X542 13313 24 446 25 CLKBUFX2 $T=1387360 1369810 0 0 $X=1387358 $Y=1369558
X543 431 24 451 25 CLKBUFX2 $T=1392880 1355050 1 0 $X=1392878 $Y=1351110
X544 13590 24 13298 25 CLKBUFX2 $T=1398860 1532170 0 0 $X=1398858 $Y=1531918
X545 13434 24 458 25 CLKBUFX2 $T=1399780 1362430 0 0 $X=1399778 $Y=1362178
X546 13590 24 13294 25 CLKBUFX2 $T=1399780 1510030 1 0 $X=1399778 $Y=1506090
X547 13659 24 366 25 CLKBUFX2 $T=1401160 1384570 1 0 $X=1401158 $Y=1380630
X548 13704 24 13272 25 CLKBUFX2 $T=1407600 1436230 1 0 $X=1407598 $Y=1432290
X549 13517 24 468 25 CLKBUFX2 $T=1415880 1369810 0 0 $X=1415878 $Y=1369558
X550 464 24 474 25 CLKBUFX2 $T=1423240 1355050 1 0 $X=1423238 $Y=1351110
X551 13723 24 473 25 CLKBUFX2 $T=1424160 1362430 0 0 $X=1424158 $Y=1362178
X552 13789 24 448 25 CLKBUFX2 $T=1430600 1502650 0 0 $X=1430598 $Y=1502398
X553 486 24 13826 25 CLKBUFX2 $T=1435660 1355050 1 0 $X=1435658 $Y=1351110
X554 398 24 12811 25 CLKBUFX2 $T=1435660 1502650 1 0 $X=1435658 $Y=1498710
X555 13948 24 13789 25 CLKBUFX2 $T=1436580 1532170 1 0 $X=1436578 $Y=1528230
X556 13928 24 13704 25 CLKBUFX2 $T=1441180 1458370 1 0 $X=1441178 $Y=1454430
X557 13928 24 13659 25 CLKBUFX2 $T=1451760 1391950 1 0 $X=1451758 $Y=1388010
X558 492 24 367 25 CLKBUFX2 $T=1454060 1355050 1 0 $X=1454058 $Y=1351110
X559 485 24 12802 25 CLKBUFX2 $T=1454520 1443610 0 0 $X=1454518 $Y=1443358
X560 457 24 516 25 CLKBUFX2 $T=1471080 1391950 0 0 $X=1471078 $Y=1391698
X561 14446 24 14158 25 CLKBUFX2 $T=1486260 1473130 1 0 $X=1486258 $Y=1469190
X562 531 24 470 25 CLKBUFX2 $T=1495000 1377190 1 0 $X=1494998 $Y=1373250
X563 526 24 342 25 CLKBUFX2 $T=1495000 1384570 0 0 $X=1494998 $Y=1384318
X564 14659 24 14282 25 CLKBUFX2 $T=1506960 1421470 1 0 $X=1506958 $Y=1417530
X565 13948 24 14194 25 CLKBUFX2 $T=1508800 1539550 0 0 $X=1508798 $Y=1539298
X566 13948 24 14446 25 CLKBUFX2 $T=1512020 1532170 1 0 $X=1512018 $Y=1528230
X567 524 24 14228 25 CLKBUFX2 $T=1515240 1428850 1 0 $X=1515238 $Y=1424910
X568 13590 24 14657 25 CLKBUFX2 $T=1517540 1539550 1 0 $X=1517538 $Y=1535610
X569 14770 24 531 25 CLKBUFX2 $T=1525360 1391950 1 0 $X=1525358 $Y=1388010
X570 14859 24 556 25 CLKBUFX2 $T=1540540 1362430 1 0 $X=1540538 $Y=1358490
X571 568 24 14659 25 CLKBUFX2 $T=1551580 1421470 0 0 $X=1551578 $Y=1421218
X572 14659 24 565 25 CLKBUFX2 $T=1563540 1384570 0 0 $X=1563538 $Y=1384318
X573 587 24 606 25 CLKBUFX2 $T=1591600 1355050 1 0 $X=1591598 $Y=1351110
X574 73 10033 49 24 25 61 MX2XL $T=1115040 1355050 0 180 $X=1111360 $Y=1351110
X575 73 10137 34 24 25 10072 MX2XL $T=1124240 1362430 0 180 $X=1120560 $Y=1358490
X576 9920 90 10343 24 25 10337 MX2XL $T=1138960 1443610 0 0 $X=1138958 $Y=1443358
X577 92 10522 10474 24 25 10657 MX2XL $T=1162420 1443610 1 0 $X=1162418 $Y=1439670
X578 92 10582 10369 24 25 10677 MX2XL $T=1162420 1465750 1 0 $X=1162418 $Y=1461810
X579 92 10645 10568 24 25 10535 MX2XL $T=1167480 1450990 1 180 $X=1163800 $Y=1450738
X580 10760 10728 10661 24 25 10508 MX2XL $T=1174380 1399330 1 180 $X=1170700 $Y=1399078
X581 92 10816 10488 24 25 10711 MX2XL $T=1184040 1458370 1 180 $X=1180360 $Y=1458118
X582 10760 11965 12026 24 25 11927 MX2XL $T=1259020 1428850 0 0 $X=1259018 $Y=1428598
X583 10760 12334 12187 24 25 12182 MX2XL $T=1283400 1443610 1 0 $X=1283398 $Y=1439670
X584 574 576 15155 24 25 15246 MX2XL $T=1559400 1369810 1 0 $X=1559398 $Y=1365870
X585 574 581 15188 24 25 15077 MX2XL $T=1563540 1355050 0 180 $X=1559860 $Y=1351110
X586 574 584 15046 24 25 15151 MX2XL $T=1564920 1362430 1 180 $X=1561240 $Y=1362178
X587 574 582 15234 24 25 15282 MX2XL $T=1562620 1355050 0 0 $X=1562618 $Y=1354798
X588 574 588 15283 24 25 15254 MX2XL $T=1573660 1362430 1 180 $X=1569980 $Y=1362178
X589 574 591 15286 24 25 15349 MX2XL $T=1575500 1355050 1 0 $X=1575498 $Y=1351110
X590 9832 9920 9825 9817 24 25 MXI2X1 $T=1098020 1436230 1 180 $X=1094800 $Y=1435978
X591 9838 9920 9944 9948 24 25 MXI2X1 $T=1102620 1377190 1 0 $X=1102618 $Y=1373250
X592 9803 9920 9909 9940 24 25 MXI2X1 $T=1104000 1384570 1 0 $X=1103998 $Y=1380630
X593 10136 9920 10051 10186 24 25 MXI2X1 $T=1127000 1450990 1 0 $X=1126998 $Y=1447050
X594 10142 9920 10240 10245 24 25 MXI2X1 $T=1130680 1414090 1 0 $X=1130678 $Y=1410150
X595 10059 92 10259 10243 24 25 MXI2X1 $T=1132060 1458370 1 0 $X=1132058 $Y=1454430
X596 10028 102 10130 10333 24 25 MXI2X1 $T=1138040 1384570 1 0 $X=1138038 $Y=1380630
X597 9949 92 10147 10338 24 25 MXI2X1 $T=1138500 1458370 1 0 $X=1138498 $Y=1454430
X598 10171 9920 10258 10297 24 25 MXI2X1 $T=1139420 1406710 1 0 $X=1139418 $Y=1402770
X599 10233 102 10296 109 24 25 MXI2X1 $T=1143100 1377190 1 0 $X=1143098 $Y=1373250
X600 10253 9920 10167 10378 24 25 MXI2X1 $T=1143560 1399330 1 0 $X=1143558 $Y=1395390
X601 10372 92 10360 10273 24 25 MXI2X1 $T=1147240 1391950 0 180 $X=1144020 $Y=1388010
X602 10165 9920 10252 10391 24 25 MXI2X1 $T=1144480 1384570 0 0 $X=1144478 $Y=1384318
X603 10358 92 10480 10271 24 25 MXI2X1 $T=1145860 1458370 1 0 $X=1145858 $Y=1454430
X604 10397 92 10383 10185 24 25 MXI2X1 $T=1149540 1377190 0 180 $X=1146320 $Y=1373250
X605 10398 92 10384 10117 24 25 MXI2X1 $T=1149540 1384570 0 180 $X=1146320 $Y=1380630
X606 10484 92 10445 10265 24 25 MXI2X1 $T=1155520 1391950 1 180 $X=1152300 $Y=1391698
X607 10392 92 10533 10501 24 25 MXI2X1 $T=1154140 1399330 0 0 $X=1154138 $Y=1399078
X608 10288 92 10500 10353 24 25 MXI2X1 $T=1154600 1458370 1 0 $X=1154598 $Y=1454430
X609 10363 102 10479 10382 24 25 MXI2X1 $T=1156440 1369810 0 0 $X=1156438 $Y=1369558
X610 12067 10760 11897 220 24 25 MXI2X1 $T=1265460 1406710 1 0 $X=1265458 $Y=1402770
X611 12216 11105 12085 11662 24 25 MXI2X1 $T=1275120 1421470 0 0 $X=1275118 $Y=1421218
X612 12341 10760 12204 11498 24 25 MXI2X1 $T=1283400 1406710 1 0 $X=1283398 $Y=1402770
X613 301 12489 12395 12513 24 25 MXI2X1 $T=1293980 1532170 0 0 $X=1293978 $Y=1531918
X614 274 12525 12522 12515 24 25 MXI2X1 $T=1301340 1443610 1 180 $X=1298120 $Y=1443358
X615 305 12489 12623 12590 24 25 MXI2X1 $T=1299500 1473130 0 0 $X=1299498 $Y=1472878
X616 308 12528 12576 12606 24 25 MXI2X1 $T=1299960 1532170 0 0 $X=1299958 $Y=1531918
X617 284 12525 12596 12593 24 25 MXI2X1 $T=1299960 1546930 0 0 $X=1299958 $Y=1546678
X618 299 12525 12571 12603 24 25 MXI2X1 $T=1300420 1421470 0 0 $X=1300418 $Y=1421218
X619 301 12528 12575 12618 24 25 MXI2X1 $T=1300880 1524790 1 0 $X=1300878 $Y=1520850
X620 308 12525 12619 12526 24 25 MXI2X1 $T=1300880 1546930 1 0 $X=1300878 $Y=1542990
X621 312 12528 12579 12227 24 25 MXI2X1 $T=1301340 1450990 0 0 $X=1301338 $Y=1450738
X622 310 12489 12563 12601 24 25 MXI2X1 $T=1302260 1414090 1 0 $X=1302258 $Y=1410150
X623 300 12528 12610 12599 24 25 MXI2X1 $T=1309620 1473130 0 180 $X=1306400 $Y=1469190
X624 310 12525 12625 12672 24 25 MXI2X1 $T=1308240 1414090 1 0 $X=1308238 $Y=1410150
X625 298 12525 12612 11806 24 25 MXI2X1 $T=1313300 1495270 0 180 $X=1310080 $Y=1491330
X626 313 12525 12640 12642 24 25 MXI2X1 $T=1313300 1517410 1 180 $X=1310080 $Y=1517158
X627 295 329 12607 12391 24 25 MXI2X1 $T=1313760 1369810 1 180 $X=1310540 $Y=1369558
X628 313 12528 12605 12637 24 25 MXI2X1 $T=1313760 1510030 0 180 $X=1310540 $Y=1506090
X629 284 12489 12639 12611 24 25 MXI2X1 $T=1311000 1539550 1 0 $X=1310998 $Y=1535610
X630 310 12675 12674 12562 24 25 MXI2X1 $T=1314220 1399330 1 180 $X=1311000 $Y=1399078
X631 300 12489 12638 12629 24 25 MXI2X1 $T=1315140 1473130 0 180 $X=1311920 $Y=1469190
X632 295 333 12705 12696 24 25 MXI2X1 $T=1319740 1369810 1 180 $X=1316520 $Y=1369558
X633 311 12525 12700 12774 24 25 MXI2X1 $T=1316980 1391950 0 0 $X=1316978 $Y=1391698
X634 309 12726 12841 12830 24 25 MXI2X1 $T=1316980 1428850 0 0 $X=1316978 $Y=1428598
X635 311 12489 12785 12780 24 25 MXI2X1 $T=1317440 1399330 1 0 $X=1317438 $Y=1395390
X636 309 12525 12775 12737 24 25 MXI2X1 $T=1317900 1414090 0 0 $X=1317898 $Y=1413838
X637 312 12525 12746 12617 24 25 MXI2X1 $T=1317900 1450990 0 0 $X=1317898 $Y=1450738
X638 305 12528 12743 12776 24 25 MXI2X1 $T=1317900 1480510 1 0 $X=1317898 $Y=1476570
X639 274 12489 12620 12702 24 25 MXI2X1 $T=1321120 1443610 1 180 $X=1317900 $Y=1443358
X640 301 12525 12713 12633 24 25 MXI2X1 $T=1321120 1510030 0 180 $X=1317900 $Y=1506090
X641 280 333 12716 331 24 25 MXI2X1 $T=1321580 1355050 1 180 $X=1318360 $Y=1354798
X642 274 12528 12826 12777 24 25 MXI2X1 $T=1319280 1436230 0 0 $X=1319278 $Y=1435978
X643 300 12726 12794 12630 24 25 MXI2X1 $T=1319280 1473130 1 0 $X=1319278 $Y=1469190
X644 298 12489 12631 12591 24 25 MXI2X1 $T=1322500 1487890 0 180 $X=1319280 $Y=1483950
X645 301 12726 12722 12738 24 25 MXI2X1 $T=1322960 1554310 0 180 $X=1319740 $Y=1550370
X646 295 341 12744 12699 24 25 MXI2X1 $T=1323420 1369810 1 180 $X=1320200 $Y=1369558
X647 300 12806 12831 12877 24 25 MXI2X1 $T=1322500 1465750 0 0 $X=1322498 $Y=1465498
X648 300 12675 12906 12907 24 25 MXI2X1 $T=1323880 1465750 1 0 $X=1323878 $Y=1461810
X649 309 12675 12803 12627 24 25 MXI2X1 $T=1327100 1421470 1 180 $X=1323880 $Y=1421218
X650 309 12528 12800 12796 24 25 MXI2X1 $T=1328020 1436230 0 0 $X=1328018 $Y=1435978
X651 298 12528 12843 12604 24 25 MXI2X1 $T=1332620 1495270 1 180 $X=1329400 $Y=1495018
X652 284 12726 12881 12795 24 25 MXI2X1 $T=1335840 1554310 0 180 $X=1332620 $Y=1550370
X653 295 355 12910 12924 24 25 MXI2X1 $T=1334000 1369810 1 0 $X=1333998 $Y=1365870
X654 313 12874 12809 12896 24 25 MXI2X1 $T=1337220 1524790 1 180 $X=1334000 $Y=1524538
X655 300 12874 12911 12842 24 25 MXI2X1 $T=1334460 1487890 1 0 $X=1334458 $Y=1483950
X656 298 12806 12888 12904 24 25 MXI2X1 $T=1337680 1502650 0 180 $X=1334460 $Y=1498710
X657 312 12675 12936 12930 24 25 MXI2X1 $T=1334920 1458370 0 0 $X=1334918 $Y=1458118
X658 308 12806 12879 12799 24 25 MXI2X1 $T=1335380 1539550 0 0 $X=1335378 $Y=1539298
X659 313 12806 12909 12781 24 25 MXI2X1 $T=1338600 1517410 0 180 $X=1335380 $Y=1513470
X660 308 12874 12940 12945 24 25 MXI2X1 $T=1335840 1554310 1 0 $X=1335838 $Y=1550370
X661 305 12806 12844 12886 24 25 MXI2X1 $T=1339060 1495270 0 180 $X=1335840 $Y=1491330
X662 313 12726 12789 12686 24 25 MXI2X1 $T=1339980 1510030 0 180 $X=1336760 $Y=1506090
X663 301 12806 12804 12801 24 25 MXI2X1 $T=1339980 1532170 0 180 $X=1336760 $Y=1528230
X664 280 368 376 377 24 25 MXI2X1 $T=1337220 1355050 1 0 $X=1337218 $Y=1351110
X665 295 369 12965 12947 24 25 MXI2X1 $T=1337220 1369810 1 0 $X=1337218 $Y=1365870
X666 305 12874 13019 13013 24 25 MXI2X1 $T=1338600 1487890 1 0 $X=1338598 $Y=1483950
X667 310 12806 12921 12836 24 25 MXI2X1 $T=1343200 1414090 0 180 $X=1339980 $Y=1410150
X668 305 12675 12972 12951 24 25 MXI2X1 $T=1343660 1473130 1 180 $X=1340440 $Y=1472878
X669 298 12874 12895 12883 24 25 MXI2X1 $T=1344120 1495270 0 180 $X=1340900 $Y=1491330
X670 310 12874 13020 12954 24 25 MXI2X1 $T=1342280 1406710 1 0 $X=1342278 $Y=1402770
X671 284 12675 13029 12956 24 25 MXI2X1 $T=1347800 1561690 0 180 $X=1344580 $Y=1557750
X672 311 12874 12920 12953 24 25 MXI2X1 $T=1348260 1391950 0 180 $X=1345040 $Y=1388010
X673 298 12675 12914 12937 24 25 MXI2X1 $T=1348260 1510030 0 180 $X=1345040 $Y=1506090
X674 301 12874 12941 12961 24 25 MXI2X1 $T=1348260 1532170 0 180 $X=1345040 $Y=1528230
X675 299 12874 12963 13035 24 25 MXI2X1 $T=1349180 1414090 0 180 $X=1345960 $Y=1410150
X676 284 12806 12967 13061 24 25 MXI2X1 $T=1346420 1532170 0 0 $X=1346418 $Y=1531918
X677 295 368 13039 12835 24 25 MXI2X1 $T=1349640 1377190 0 180 $X=1346420 $Y=1373250
X678 298 12726 13041 12898 24 25 MXI2X1 $T=1349640 1495270 0 180 $X=1346420 $Y=1491330
X679 280 369 12968 13064 24 25 MXI2X1 $T=1347340 1362430 1 0 $X=1347338 $Y=1358490
X680 309 12874 13045 12949 24 25 MXI2X1 $T=1350560 1436230 0 180 $X=1347340 $Y=1432290
X681 13057 44 389 13104 24 25 MXI2X1 $T=1349180 1384570 0 0 $X=1349178 $Y=1384318
X682 299 12675 13093 13108 24 25 MXI2X1 $T=1349180 1428850 1 0 $X=1349178 $Y=1424910
X683 311 12806 13067 13030 24 25 MXI2X1 $T=1352860 1377190 0 180 $X=1349640 $Y=1373250
X684 295 371 13136 13117 24 25 MXI2X1 $T=1351480 1362430 0 0 $X=1351478 $Y=1362178
X685 308 12675 13134 13139 24 25 MXI2X1 $T=1351480 1561690 0 0 $X=1351478 $Y=1561438
X686 312 12874 13138 13149 24 25 MXI2X1 $T=1352400 1465750 1 0 $X=1352398 $Y=1461810
X687 313 12675 13167 13065 24 25 MXI2X1 $T=1352400 1510030 0 0 $X=1352398 $Y=1509778
X688 311 12675 12962 13056 24 25 MXI2X1 $T=1355620 1391950 0 180 $X=1352400 $Y=1388010
X689 308 12726 13123 13146 24 25 MXI2X1 $T=1352860 1554310 1 0 $X=1352858 $Y=1550370
X690 13122 74 12245 13150 24 25 MXI2X1 $T=1353320 1487890 0 0 $X=1353318 $Y=1487638
X691 312 12726 13125 12827 24 25 MXI2X1 $T=1356540 1473130 0 180 $X=1353320 $Y=1469190
X692 274 12675 13182 13027 24 25 MXI2X1 $T=1353780 1436230 0 0 $X=1353778 $Y=1435978
X693 301 12675 13112 13186 24 25 MXI2X1 $T=1353780 1524790 1 0 $X=1353778 $Y=1520850
X694 311 12726 13126 13170 24 25 MXI2X1 $T=1354240 1391950 0 0 $X=1354238 $Y=1391698
X695 299 12726 13174 13156 24 25 MXI2X1 $T=1354240 1406710 0 0 $X=1354238 $Y=1406458
X696 280 371 13154 13240 24 25 MXI2X1 $T=1358380 1362430 1 0 $X=1358378 $Y=1358490
X697 13187 74 12021 13248 24 25 MXI2X1 $T=1359760 1495270 1 0 $X=1359758 $Y=1491330
X698 13188 74 12193 13233 24 25 MXI2X1 $T=1360680 1384570 1 0 $X=1360678 $Y=1380630
X699 13226 74 11882 13257 24 25 MXI2X1 $T=1362520 1406710 0 0 $X=1362518 $Y=1406458
X700 309 13241 13155 13258 24 25 MXI2X1 $T=1362520 1436230 0 0 $X=1362518 $Y=1435978
X701 13230 74 12081 13291 24 25 MXI2X1 $T=1362520 1524790 1 0 $X=1362518 $Y=1520850
X702 13251 417 12018 13177 24 25 MXI2X1 $T=1365740 1495270 1 180 $X=1362520 $Y=1495018
X703 13231 44 408 13284 24 25 MXI2X1 $T=1362980 1458370 1 0 $X=1362978 $Y=1454430
X704 13234 74 12237 13269 24 25 MXI2X1 $T=1363440 1399330 0 0 $X=1363438 $Y=1399078
X705 13238 74 12084 13265 24 25 MXI2X1 $T=1363440 1517410 0 0 $X=1363438 $Y=1517158
X706 13245 74 12252 13281 24 25 MXI2X1 $T=1363900 1458370 0 0 $X=1363898 $Y=1458118
X707 13247 44 12251 13286 24 25 MXI2X1 $T=1363900 1502650 1 0 $X=1363898 $Y=1498710
X708 305 12726 13261 13055 24 25 MXI2X1 $T=1364820 1473130 0 0 $X=1364818 $Y=1472878
X709 13181 414 415 13301 24 25 MXI2X1 $T=1367120 1391950 1 0 $X=1367118 $Y=1388010
X710 311 13312 13311 13367 24 25 MXI2X1 $T=1368960 1399330 1 0 $X=1368958 $Y=1395390
X711 309 13313 13356 13362 24 25 MXI2X1 $T=1368960 1414090 0 0 $X=1368958 $Y=1413838
X712 13295 44 422 13363 24 25 MXI2X1 $T=1368960 1436230 1 0 $X=1368958 $Y=1432290
X713 313 13241 13365 13292 24 25 MXI2X1 $T=1368960 1524790 1 0 $X=1368958 $Y=1520850
X714 310 13241 13361 13474 24 25 MXI2X1 $T=1369880 1414090 1 0 $X=1369878 $Y=1410150
X715 301 13312 13354 13376 24 25 MXI2X1 $T=1370340 1532170 1 0 $X=1370338 $Y=1528230
X716 295 411 13319 13137 24 25 MXI2X1 $T=1373560 1377190 0 180 $X=1370340 $Y=1373250
X717 13306 413 426 13394 24 25 MXI2X1 $T=1370800 1369810 1 0 $X=1370798 $Y=1365870
X718 299 13313 13381 13385 24 25 MXI2X1 $T=1370800 1421470 0 0 $X=1370798 $Y=1421218
X719 13349 74 12351 13403 24 25 MXI2X1 $T=1371260 1436230 0 0 $X=1371258 $Y=1435978
X720 13276 74 12020 13386 24 25 MXI2X1 $T=1371260 1473130 0 0 $X=1371258 $Y=1472878
X721 305 13313 13303 13419 24 25 MXI2X1 $T=1371260 1495270 0 0 $X=1371258 $Y=1495018
X722 301 13313 13266 13014 24 25 MXI2X1 $T=1374480 1546930 1 180 $X=1371260 $Y=1546678
X723 280 411 429 430 24 25 MXI2X1 $T=1372180 1355050 1 0 $X=1372178 $Y=1351110
X724 301 13434 13287 13173 24 25 MXI2X1 $T=1375400 1524790 1 180 $X=1372180 $Y=1524538
X725 13371 74 11947 13400 24 25 MXI2X1 $T=1372640 1443610 1 0 $X=1372638 $Y=1439670
X726 284 13312 13399 13409 24 25 MXI2X1 $T=1373560 1532170 1 0 $X=1373558 $Y=1528230
X727 301 13241 13160 13279 24 25 MXI2X1 $T=1378620 1554310 1 180 $X=1375400 $Y=1554058
X728 280 423 13414 13380 24 25 MXI2X1 $T=1375860 1355050 1 0 $X=1375858 $Y=1351110
X729 309 13312 13412 13307 24 25 MXI2X1 $T=1379540 1399330 0 180 $X=1376320 $Y=1395390
X730 295 423 13388 13440 24 25 MXI2X1 $T=1377240 1362430 1 0 $X=1377238 $Y=1358490
X731 300 13434 13423 13350 24 25 MXI2X1 $T=1381380 1458370 0 180 $X=1378160 $Y=1454430
X732 305 13241 13431 13387 24 25 MXI2X1 $T=1379080 1495270 0 0 $X=1379078 $Y=1495018
X733 309 13434 13472 13369 24 25 MXI2X1 $T=1379540 1436230 0 0 $X=1379538 $Y=1435978
X734 284 13241 13435 13355 24 25 MXI2X1 $T=1379540 1561690 1 0 $X=1379538 $Y=1557750
X735 284 13313 13428 13270 24 25 MXI2X1 $T=1382760 1546930 1 180 $X=1379540 $Y=1546678
X736 300 13241 13441 13420 24 25 MXI2X1 $T=1380000 1480510 1 0 $X=1379998 $Y=1476570
X737 298 13313 13439 13408 24 25 MXI2X1 $T=1384140 1510030 0 180 $X=1380920 $Y=1506090
X738 274 13241 13364 13437 24 25 MXI2X1 $T=1385060 1458370 0 180 $X=1381840 $Y=1454430
X739 311 13241 13529 13477 24 25 MXI2X1 $T=1382760 1399330 1 0 $X=1382758 $Y=1395390
X740 311 13313 13389 13436 24 25 MXI2X1 $T=1388740 1377190 1 180 $X=1385520 $Y=1376938
X741 310 13434 13508 13525 24 25 MXI2X1 $T=1385980 1406710 0 0 $X=1385978 $Y=1406458
X742 274 13434 13493 13357 24 25 MXI2X1 $T=1385980 1450990 1 0 $X=1385978 $Y=1447050
X743 284 13434 13500 13483 24 25 MXI2X1 $T=1389200 1524790 1 180 $X=1385980 $Y=1524538
X744 300 13312 13504 13418 24 25 MXI2X1 $T=1389660 1480510 0 180 $X=1386440 $Y=1476570
X745 312 13434 13515 13532 24 25 MXI2X1 $T=1386900 1450990 0 0 $X=1386898 $Y=1450738
X746 312 13313 13486 13533 24 25 MXI2X1 $T=1386900 1458370 0 0 $X=1386898 $Y=1458118
X747 312 13241 13495 13512 24 25 MXI2X1 $T=1386900 1465750 0 0 $X=1386898 $Y=1465498
X748 305 13312 13498 13411 24 25 MXI2X1 $T=1390120 1487890 0 180 $X=1386900 $Y=1483950
X749 298 13241 13442 13366 24 25 MXI2X1 $T=1390120 1510030 1 180 $X=1386900 $Y=1509778
X750 313 13517 13583 13582 24 25 MXI2X1 $T=1387360 1517410 0 0 $X=1387358 $Y=1517158
X751 310 13312 13538 13481 24 25 MXI2X1 $T=1388280 1414090 1 0 $X=1388278 $Y=1410150
X752 305 13434 13574 13479 24 25 MXI2X1 $T=1388280 1495270 1 0 $X=1388278 $Y=1491330
X753 298 13434 13597 13513 24 25 MXI2X1 $T=1388280 1502650 0 0 $X=1388278 $Y=1502398
X754 274 13313 13478 13382 24 25 MXI2X1 $T=1391500 1436230 1 180 $X=1388280 $Y=1435978
X755 313 13313 13494 13406 24 25 MXI2X1 $T=1391500 1524790 0 180 $X=1388280 $Y=1520850
X756 308 13434 13518 13510 24 25 MXI2X1 $T=1391500 1539550 0 180 $X=1388280 $Y=1535610
X757 295 438 13521 437 24 25 MXI2X1 $T=1391960 1362430 1 180 $X=1388740 $Y=1362178
X758 295 439 13579 13509 24 25 MXI2X1 $T=1389200 1369810 0 0 $X=1389198 $Y=1369558
X759 308 13241 13506 13575 24 25 MXI2X1 $T=1389660 1554310 0 0 $X=1389658 $Y=1554058
X760 299 13241 13531 13496 24 25 MXI2X1 $T=1393800 1428850 1 180 $X=1390580 $Y=1428598
X761 299 450 13581 13585 24 25 MXI2X1 $T=1391500 1428850 1 0 $X=1391498 $Y=1424910
X762 280 439 13615 13516 24 25 MXI2X1 $T=1391960 1355050 0 0 $X=1391958 $Y=1354798
X763 295 452 13573 13610 24 25 MXI2X1 $T=1392880 1384570 1 0 $X=1392878 $Y=1380630
X764 308 13313 13594 13514 24 25 MXI2X1 $T=1392880 1546930 0 0 $X=1392878 $Y=1546678
X765 311 13434 13605 13580 24 25 MXI2X1 $T=1399780 1384570 1 180 $X=1396560 $Y=1384318
X766 274 13312 13587 13491 24 25 MXI2X1 $T=1399780 1436230 1 180 $X=1396560 $Y=1435978
X767 299 13434 13619 13526 24 25 MXI2X1 $T=1397020 1414090 1 0 $X=1397018 $Y=1410150
X768 305 13517 13596 13678 24 25 MXI2X1 $T=1397020 1495270 1 0 $X=1397018 $Y=1491330
X769 274 450 13607 13523 24 25 MXI2X1 $T=1400240 1428850 1 180 $X=1397020 $Y=1428598
X770 298 13312 13601 13499 24 25 MXI2X1 $T=1400240 1502650 1 180 $X=1397020 $Y=1502398
X771 313 13312 13611 13536 24 25 MXI2X1 $T=1400240 1524790 0 180 $X=1397020 $Y=1520850
X772 308 13312 13612 13519 24 25 MXI2X1 $T=1400240 1539550 0 180 $X=1397020 $Y=1535610
X773 280 452 13598 456 24 25 MXI2X1 $T=1401620 1355050 1 180 $X=1398400 $Y=1354798
X774 312 13312 13622 13593 24 25 MXI2X1 $T=1401620 1458370 0 180 $X=1398400 $Y=1454430
X775 313 13434 13603 13502 24 25 MXI2X1 $T=1402540 1517410 0 180 $X=1399320 $Y=1513470
X776 299 13312 13599 13501 24 25 MXI2X1 $T=1403000 1421470 1 180 $X=1399780 $Y=1421218
X777 300 13517 13650 13492 24 25 MXI2X1 $T=1404380 1473130 1 180 $X=1401160 $Y=1472878
X778 309 13517 13674 13689 24 25 MXI2X1 $T=1402540 1428850 0 0 $X=1402538 $Y=1428598
X779 310 13517 13681 13697 24 25 MXI2X1 $T=1403460 1391950 0 0 $X=1403458 $Y=1391698
X780 305 450 13684 13672 24 25 MXI2X1 $T=1403460 1487890 1 0 $X=1403458 $Y=1483950
X781 313 450 13685 13699 24 25 MXI2X1 $T=1403460 1524790 1 0 $X=1403458 $Y=1520850
X782 308 13517 13675 13606 24 25 MXI2X1 $T=1406680 1532170 0 180 $X=1403460 $Y=1528230
X783 310 450 13693 13707 24 25 MXI2X1 $T=1404380 1406710 0 0 $X=1404378 $Y=1406458
X784 274 13517 13719 13661 24 25 MXI2X1 $T=1404380 1458370 1 0 $X=1404378 $Y=1454430
X785 295 462 13591 13592 24 25 MXI2X1 $T=1407600 1362430 1 180 $X=1404380 $Y=1362178
X786 295 463 13686 13537 24 25 MXI2X1 $T=1408060 1384570 0 180 $X=1404840 $Y=1380630
X787 310 464 13687 13673 24 25 MXI2X1 $T=1408060 1399330 1 180 $X=1404840 $Y=1399078
X788 300 450 13539 13654 24 25 MXI2X1 $T=1408060 1473130 1 180 $X=1404840 $Y=1472878
X789 308 464 13692 13679 24 25 MXI2X1 $T=1408520 1546930 1 180 $X=1405300 $Y=1546678
X790 308 450 13578 13616 24 25 MXI2X1 $T=1408980 1554310 1 180 $X=1405760 $Y=1554058
X791 298 450 13705 13721 24 25 MXI2X1 $T=1406220 1495270 0 0 $X=1406218 $Y=1495018
X792 298 13517 13682 13759 24 25 MXI2X1 $T=1406220 1502650 0 0 $X=1406218 $Y=1502398
X793 274 464 13653 13694 24 25 MXI2X1 $T=1409440 1443610 0 180 $X=1406220 $Y=1439670
X794 312 450 13720 13712 24 25 MXI2X1 $T=1406680 1465750 1 0 $X=1406678 $Y=1461810
X795 301 13517 13708 13724 24 25 MXI2X1 $T=1407140 1532170 1 0 $X=1407138 $Y=1528230
X796 280 463 13706 13695 24 25 MXI2X1 $T=1410360 1355050 0 180 $X=1407140 $Y=1351110
X797 311 13517 13666 13715 24 25 MXI2X1 $T=1408520 1391950 1 0 $X=1408518 $Y=1388010
X798 311 462 13700 13765 24 25 MXI2X1 $T=1410820 1362430 0 0 $X=1410818 $Y=1362178
X799 305 461 13755 13669 24 25 MXI2X1 $T=1411740 1480510 1 0 $X=1411738 $Y=1476570
X800 274 461 13751 13703 24 25 MXI2X1 $T=1415420 1450990 0 180 $X=1412200 $Y=1447050
X801 300 464 13769 13683 24 25 MXI2X1 $T=1417260 1465750 0 180 $X=1414040 $Y=1461810
X802 301 450 13691 13764 24 25 MXI2X1 $T=1417260 1554310 1 180 $X=1414040 $Y=1554058
X803 284 13517 13667 13752 24 25 MXI2X1 $T=1418640 1539550 0 180 $X=1415420 $Y=1535610
X804 311 450 13776 13677 24 25 MXI2X1 $T=1419560 1399330 0 180 $X=1416340 $Y=1395390
X805 299 13517 13709 13777 24 25 MXI2X1 $T=1420020 1414090 0 180 $X=1416800 $Y=1410150
X806 313 461 13757 13676 24 25 MXI2X1 $T=1420480 1517410 0 180 $X=1417260 $Y=1513470
X807 305 13826 13828 13840 24 25 MXI2X1 $T=1420020 1480510 0 0 $X=1420018 $Y=1480258
X808 284 450 13846 13842 24 25 MXI2X1 $T=1420480 1554310 1 0 $X=1420478 $Y=1550370
X809 300 461 13781 13713 24 25 MXI2X1 $T=1423700 1473130 0 180 $X=1420480 $Y=1469190
X810 471 464 13825 13773 24 25 MXI2X1 $T=1424160 1362430 0 180 $X=1420940 $Y=1358490
X811 311 13826 13838 13862 24 25 MXI2X1 $T=1421400 1391950 0 0 $X=1421398 $Y=1391698
X812 309 461 13796 13868 24 25 MXI2X1 $T=1421400 1421470 0 0 $X=1421398 $Y=1421218
X813 298 13826 13863 13881 24 25 MXI2X1 $T=1421400 1510030 1 0 $X=1421398 $Y=1506090
X814 472 464 13760 13663 24 25 MXI2X1 $T=1424620 1369810 1 180 $X=1421400 $Y=1369558
X815 311 464 13722 13788 24 25 MXI2X1 $T=1424620 1377190 1 180 $X=1421400 $Y=1376938
X816 13844 464 13790 13690 24 25 MXI2X1 $T=1424620 1421470 0 180 $X=1421400 $Y=1417530
X817 305 464 13782 13534 24 25 MXI2X1 $T=1424620 1487890 1 180 $X=1421400 $Y=1487638
X818 313 464 13783 13711 24 25 MXI2X1 $T=1424620 1517410 0 180 $X=1421400 $Y=1513470
X819 298 461 13884 13792 24 25 MXI2X1 $T=1421860 1502650 1 0 $X=1421858 $Y=1498710
X820 309 450 13829 13750 24 25 MXI2X1 $T=1425080 1428850 1 180 $X=1421860 $Y=1428598
X821 13850 464 13835 13833 24 25 MXI2X1 $T=1425540 1399330 1 180 $X=1422320 $Y=1399078
X822 301 461 13843 13837 24 25 MXI2X1 $T=1426000 1524790 0 180 $X=1422780 $Y=1520850
X823 308 461 13763 13680 24 25 MXI2X1 $T=1426000 1546930 1 180 $X=1422780 $Y=1546678
X824 274 13826 13855 13832 24 25 MXI2X1 $T=1423240 1443610 1 0 $X=1423238 $Y=1439670
X825 312 464 13897 13830 24 25 MXI2X1 $T=1424160 1458370 1 0 $X=1424158 $Y=1454430
X826 295 476 13880 13893 24 25 MXI2X1 $T=1426000 1362430 1 0 $X=1425998 $Y=1358490
X827 13836 13885 13879 13851 24 25 MXI2X1 $T=1429680 1443610 1 180 $X=1426460 $Y=1443358
X828 298 464 13883 13834 24 25 MXI2X1 $T=1430600 1487890 1 180 $X=1427380 $Y=1487638
X829 13891 13932 13859 13882 24 25 MXI2X1 $T=1431060 1377190 1 180 $X=1427840 $Y=1376938
X830 13891 13885 13878 13784 24 25 MXI2X1 $T=1431060 1391950 1 180 $X=1427840 $Y=1391698
X831 299 13826 13874 13839 24 25 MXI2X1 $T=1429680 1414090 0 0 $X=1429678 $Y=1413838
X832 310 461 13898 13827 24 25 MXI2X1 $T=1431060 1406710 0 0 $X=1431058 $Y=1406458
X833 284 461 13936 13866 24 25 MXI2X1 $T=1431520 1546930 0 0 $X=1431518 $Y=1546678
X834 13894 13885 13926 13857 24 25 MXI2X1 $T=1434740 1524790 0 180 $X=1431520 $Y=1520850
X835 472 483 13931 13858 24 25 MXI2X1 $T=1436120 1369810 1 180 $X=1432900 $Y=1369558
X836 13877 13885 13841 13824 24 25 MXI2X1 $T=1436120 1487890 1 180 $X=1432900 $Y=1487638
X837 13891 13980 13869 13873 24 25 MXI2X1 $T=1437040 1391950 1 180 $X=1433820 $Y=1391698
X838 13877 13932 13934 13860 24 25 MXI2X1 $T=1437500 1458370 1 180 $X=1434280 $Y=1458118
X839 13877 13980 13942 13875 24 25 MXI2X1 $T=1440260 1480510 0 180 $X=1437040 $Y=1476570
X840 284 464 13943 13872 24 25 MXI2X1 $T=1437500 1539550 0 0 $X=1437498 $Y=1539298
X841 13836 13959 13977 13992 24 25 MXI2X1 $T=1437960 1458370 1 0 $X=1437958 $Y=1454430
X842 13877 13959 14003 13995 24 25 MXI2X1 $T=1437960 1487890 0 0 $X=1437958 $Y=1487638
X843 13844 13996 13963 13957 24 25 MXI2X1 $T=1441180 1436230 0 180 $X=1437960 $Y=1432290
X844 13894 13996 13967 13887 24 25 MXI2X1 $T=1441180 1510030 1 180 $X=1437960 $Y=1509778
X845 13894 13932 13938 13870 24 25 MXI2X1 $T=1441180 1524790 1 180 $X=1437960 $Y=1524538
X846 284 13826 14004 14047 24 25 MXI2X1 $T=1438880 1546930 0 0 $X=1438878 $Y=1546678
X847 13894 13959 13956 13972 24 25 MXI2X1 $T=1442100 1524790 0 180 $X=1438880 $Y=1520850
X848 13836 13932 13979 14061 24 25 MXI2X1 $T=1439340 1450990 0 0 $X=1439338 $Y=1450738
X849 472 489 13981 13961 24 25 MXI2X1 $T=1442560 1377190 0 180 $X=1439340 $Y=1373250
X850 13877 13996 13974 14042 24 25 MXI2X1 $T=1440260 1480510 1 0 $X=1440258 $Y=1476570
X851 13844 13932 13991 13984 24 25 MXI2X1 $T=1443480 1428850 0 180 $X=1440260 $Y=1424910
X852 13894 13980 13944 13864 24 25 MXI2X1 $T=1443480 1532170 1 180 $X=1440260 $Y=1531918
X853 13844 13980 14034 14006 24 25 MXI2X1 $T=1440720 1406710 1 0 $X=1440718 $Y=1402770
X854 14032 13959 14048 14116 24 25 MXI2X1 $T=1441640 1510030 0 0 $X=1441638 $Y=1509778
X855 13836 13980 14035 13973 24 25 MXI2X1 $T=1444860 1436230 0 180 $X=1441640 $Y=1432290
X856 13877 14131 14036 13935 24 25 MXI2X1 $T=1444860 1465750 0 180 $X=1441640 $Y=1461810
X857 472 488 13968 13849 24 25 MXI2X1 $T=1442560 1369810 1 0 $X=1442558 $Y=1365870
X858 14032 13932 13999 13997 24 25 MXI2X1 $T=1442560 1539550 0 0 $X=1442558 $Y=1539298
X859 14032 497 14055 14037 24 25 MXI2X1 $T=1447620 1502650 1 180 $X=1444400 $Y=1502398
X860 13844 13959 14064 14119 24 25 MXI2X1 $T=1445320 1436230 1 0 $X=1445318 $Y=1432290
X861 13844 13885 14120 13966 24 25 MXI2X1 $T=1448540 1428850 1 0 $X=1448538 $Y=1424910
X862 13836 13996 14069 14049 24 25 MXI2X1 $T=1451760 1458370 1 180 $X=1448540 $Y=1458118
X863 14032 13885 14076 13990 24 25 MXI2X1 $T=1451760 1532170 1 180 $X=1448540 $Y=1531918
X864 13891 13996 14129 14041 24 25 MXI2X1 $T=1449000 1377190 1 0 $X=1448998 $Y=1373250
X865 13891 497 14045 14138 24 25 MXI2X1 $T=1449920 1406710 1 0 $X=1449918 $Y=1402770
X866 13894 497 14121 14054 24 25 MXI2X1 $T=1453140 1502650 0 180 $X=1449920 $Y=1498710
X867 13894 14131 14132 14043 24 25 MXI2X1 $T=1454060 1487890 0 180 $X=1450840 $Y=1483950
X868 13891 14168 14170 14188 24 25 MXI2X1 $T=1454980 1399330 1 0 $X=1454978 $Y=1395390
X869 14032 14168 14189 14181 24 25 MXI2X1 $T=1454980 1502650 1 0 $X=1454978 $Y=1498710
X870 308 13826 14191 14190 24 25 MXI2X1 $T=1454980 1546930 0 0 $X=1454978 $Y=1546678
X871 13891 13959 14156 14157 24 25 MXI2X1 $T=1458200 1391950 1 180 $X=1454980 $Y=1391698
X872 14032 13996 14136 14046 24 25 MXI2X1 $T=1458200 1532170 1 180 $X=1454980 $Y=1531918
X873 13844 14131 14171 14130 24 25 MXI2X1 $T=1459120 1421470 0 180 $X=1455900 $Y=1417530
X874 13836 497 14172 14265 24 25 MXI2X1 $T=1457280 1458370 0 0 $X=1457278 $Y=1458118
X875 13877 497 14143 14051 24 25 MXI2X1 $T=1460500 1480510 1 180 $X=1457280 $Y=1480258
X876 471 509 14167 14068 24 25 MXI2X1 $T=1461880 1377190 0 180 $X=1458660 $Y=1373250
X877 13891 14131 14231 14148 24 25 MXI2X1 $T=1463260 1391950 1 180 $X=1460040 $Y=1391698
X878 13877 14168 14238 14164 24 25 MXI2X1 $T=1463720 1480510 1 180 $X=1460500 $Y=1480258
X879 14032 14131 14229 14123 24 25 MXI2X1 $T=1463720 1517410 1 180 $X=1460500 $Y=1517158
X880 14230 13980 14278 14186 24 25 MXI2X1 $T=1461880 1539550 0 0 $X=1461878 $Y=1539298
X881 13894 14168 14245 14176 24 25 MXI2X1 $T=1465100 1495270 0 180 $X=1461880 $Y=1491330
X882 13836 14273 14174 14267 24 25 MXI2X1 $T=1469240 1458370 1 180 $X=1466020 $Y=1458118
X883 13844 14168 14275 14233 24 25 MXI2X1 $T=1470620 1428850 0 180 $X=1467400 $Y=1424910
X884 13894 14318 14260 14274 24 25 MXI2X1 $T=1470620 1510030 0 180 $X=1467400 $Y=1506090
X885 13877 14273 14169 14268 24 25 MXI2X1 $T=1471540 1487890 0 180 $X=1468320 $Y=1483950
X886 14032 13980 14284 14236 24 25 MXI2X1 $T=1475220 1546930 0 180 $X=1472000 $Y=1542990
X887 14230 14273 14353 14351 24 25 MXI2X1 $T=1472460 1510030 1 0 $X=1472458 $Y=1506090
X888 13844 14318 14336 14321 24 25 MXI2X1 $T=1475680 1428850 0 180 $X=1472460 $Y=1424910
X889 13844 497 14234 14317 24 25 MXI2X1 $T=1475680 1436230 0 180 $X=1472460 $Y=1432290
X890 13877 14318 14330 14249 24 25 MXI2X1 $T=1475680 1458370 1 180 $X=1472460 $Y=1458118
X891 14230 497 14322 14331 24 25 MXI2X1 $T=1475680 1480510 1 180 $X=1472460 $Y=1480258
X892 14032 14273 14277 14140 24 25 MXI2X1 $T=1475680 1532170 0 180 $X=1472460 $Y=1528230
X893 310 13826 14323 14313 24 25 MXI2X1 $T=1476140 1414090 0 180 $X=1472920 $Y=1410150
X894 14230 13996 14343 14315 24 25 MXI2X1 $T=1476600 1495270 1 180 $X=1473380 $Y=1495018
X895 13894 14358 14344 14339 24 25 MXI2X1 $T=1476600 1502650 0 180 $X=1473380 $Y=1498710
X896 14032 14358 14342 14252 24 25 MXI2X1 $T=1476600 1517410 1 180 $X=1473380 $Y=1517158
X897 471 517 14225 513 24 25 MXI2X1 $T=1477060 1355050 0 180 $X=1473840 $Y=1351110
X898 13836 14131 14283 14235 24 25 MXI2X1 $T=1477060 1443610 1 180 $X=1473840 $Y=1443358
X899 13844 14358 14346 14328 24 25 MXI2X1 $T=1477520 1414090 1 180 $X=1474300 $Y=1413838
X900 14032 14318 14341 14263 24 25 MXI2X1 $T=1477520 1510030 1 180 $X=1474300 $Y=1509778
X901 312 13826 14347 14375 24 25 MXI2X1 $T=1474760 1436230 0 0 $X=1474758 $Y=1435978
X902 300 13826 14364 14412 24 25 MXI2X1 $T=1474760 1458370 1 0 $X=1474758 $Y=1454430
X903 14230 13885 14439 14352 24 25 MXI2X1 $T=1474760 1539550 0 0 $X=1474758 $Y=1539298
X904 472 505 14261 14340 24 25 MXI2X1 $T=1477980 1377190 0 180 $X=1474760 $Y=1373250
X905 13891 14358 14350 14128 24 25 MXI2X1 $T=1477980 1384570 0 180 $X=1474760 $Y=1380630
X906 13894 14273 14333 14259 24 25 MXI2X1 $T=1477980 1480510 0 180 $X=1474760 $Y=1476570
X907 14230 14358 14372 14380 24 25 MXI2X1 $T=1476600 1510030 1 0 $X=1476598 $Y=1506090
X908 14230 13932 14360 14332 24 25 MXI2X1 $T=1479820 1532170 1 180 $X=1476600 $Y=1531918
X909 14356 13932 14320 14379 24 25 MXI2X1 $T=1482580 1414090 0 180 $X=1479360 $Y=1410150
X910 14230 14131 14365 14438 24 25 MXI2X1 $T=1482120 1487890 1 0 $X=1482118 $Y=1483950
X911 14255 13932 14368 14455 24 25 MXI2X1 $T=1482120 1524790 0 0 $X=1482118 $Y=1524538
X912 13836 14318 14419 14329 24 25 MXI2X1 $T=1485800 1458370 0 180 $X=1482580 $Y=1454430
X913 471 523 14435 14349 24 25 MXI2X1 $T=1483040 1377190 1 0 $X=1483038 $Y=1373250
X914 14421 13932 14367 14451 24 25 MXI2X1 $T=1483040 1428850 0 0 $X=1483038 $Y=1428598
X915 301 13826 14373 14443 24 25 MXI2X1 $T=1483040 1554310 1 0 $X=1483038 $Y=1550370
X916 472 515 522 518 24 25 MXI2X1 $T=1486260 1355050 0 180 $X=1483040 $Y=1351110
X917 13891 14318 14428 14355 24 25 MXI2X1 $T=1486260 1384570 0 180 $X=1483040 $Y=1380630
X918 13891 14273 14429 14345 24 25 MXI2X1 $T=1486260 1391950 0 180 $X=1483040 $Y=1388010
X919 13850 13980 14425 14319 24 25 MXI2X1 $T=1486260 1399330 0 180 $X=1483040 $Y=1395390
X920 13836 14168 14430 14361 24 25 MXI2X1 $T=1486260 1436230 1 180 $X=1483040 $Y=1435978
X921 14356 13980 14374 14449 24 25 MXI2X1 $T=1483500 1421470 1 0 $X=1483498 $Y=1417530
X922 13836 14358 14436 14371 24 25 MXI2X1 $T=1487180 1450990 1 180 $X=1483960 $Y=1450738
X923 14450 13932 14426 14166 24 25 MXI2X1 $T=1487180 1465750 1 180 $X=1483960 $Y=1465498
X924 13877 14358 14434 14348 24 25 MXI2X1 $T=1487180 1473130 1 180 $X=1483960 $Y=1472878
X925 471 520 14437 14377 24 25 MXI2X1 $T=1487640 1369810 0 180 $X=1484420 $Y=1365870
X926 13844 14273 14444 14359 24 25 MXI2X1 $T=1488560 1421470 1 180 $X=1485340 $Y=1421218
X927 14356 13996 14472 14513 24 25 MXI2X1 $T=1488560 1421470 1 0 $X=1488558 $Y=1417530
X928 14421 13885 14514 14515 24 25 MXI2X1 $T=1489020 1443610 0 0 $X=1489018 $Y=1443358
X929 14467 13996 14473 14526 24 25 MXI2X1 $T=1489480 1524790 0 0 $X=1489478 $Y=1524538
X930 13850 13932 14531 14427 24 25 MXI2X1 $T=1489940 1399330 0 0 $X=1489938 $Y=1399078
X931 14467 13932 14549 14532 24 25 MXI2X1 $T=1490400 1532170 0 0 $X=1490398 $Y=1531918
X932 472 501 14422 14334 24 25 MXI2X1 $T=1491780 1355050 1 0 $X=1491778 $Y=1351110
X933 472 509 14511 14537 24 25 MXI2X1 $T=1491780 1377190 1 0 $X=1491778 $Y=1373250
X934 14450 13996 14463 14536 24 25 MXI2X1 $T=1491780 1473130 0 0 $X=1491778 $Y=1472878
X935 14450 13885 14518 14362 24 25 MXI2X1 $T=1495000 1450990 1 180 $X=1491780 $Y=1450738
X936 14230 13959 14519 14447 24 25 MXI2X1 $T=1495000 1480510 1 180 $X=1491780 $Y=1480258
X937 14421 13996 14586 14585 24 25 MXI2X1 $T=1492240 1443610 0 0 $X=1492238 $Y=1443358
X938 14467 13980 14550 14647 24 25 MXI2X1 $T=1493620 1546930 1 0 $X=1493618 $Y=1542990
X939 472 523 14553 534 24 25 MXI2X1 $T=1494080 1355050 0 0 $X=1494078 $Y=1354798
X940 14421 13980 14556 14457 24 25 MXI2X1 $T=1498220 1428850 0 180 $X=1495000 $Y=1424910
X941 13850 13996 14548 14567 24 25 MXI2X1 $T=1495920 1384570 1 0 $X=1495918 $Y=1380630
X942 14450 497 14544 14640 24 25 MXI2X1 $T=1500520 1473130 0 0 $X=1500518 $Y=1472878
X943 14255 13996 14660 14570 24 25 MXI2X1 $T=1500520 1480510 0 0 $X=1500518 $Y=1480258
X944 472 510 535 532 24 25 MXI2X1 $T=1503740 1355050 0 180 $X=1500520 $Y=1351110
X945 14450 13980 14619 14525 24 25 MXI2X1 $T=1503740 1450990 1 180 $X=1500520 $Y=1450738
X946 14467 497 14620 14431 24 25 MXI2X1 $T=1503740 1510030 0 180 $X=1500520 $Y=1506090
X947 14230 14168 14654 14564 24 25 MXI2X1 $T=1501900 1502650 0 0 $X=1501898 $Y=1502398
X948 13850 13885 14629 14543 24 25 MXI2X1 $T=1505120 1391950 0 180 $X=1501900 $Y=1388010
X949 14255 13980 14634 14542 24 25 MXI2X1 $T=1502360 1532170 1 0 $X=1502358 $Y=1528230
X950 14356 497 14639 14551 24 25 MXI2X1 $T=1502820 1399330 1 0 $X=1502818 $Y=1395390
X951 14467 14273 14673 14676 24 25 MXI2X1 $T=1505580 1532170 1 0 $X=1505578 $Y=1528230
X952 14421 14131 14677 14670 24 25 MXI2X1 $T=1506960 1450990 1 0 $X=1506958 $Y=1447050
X953 13850 14131 14662 14638 24 25 MXI2X1 $T=1510180 1399330 0 180 $X=1506960 $Y=1395390
X954 14421 497 14555 14554 24 25 MXI2X1 $T=1510180 1428850 0 180 $X=1506960 $Y=1424910
X955 14450 14131 14762 14678 24 25 MXI2X1 $T=1507420 1465750 0 0 $X=1507418 $Y=1465498
X956 13850 13959 14685 14731 24 25 MXI2X1 $T=1507880 1399330 0 0 $X=1507878 $Y=1399078
X957 14255 13959 14740 14667 24 25 MXI2X1 $T=1508340 1487890 0 0 $X=1508338 $Y=1487638
X958 472 517 540 538 24 25 MXI2X1 $T=1508800 1355050 1 0 $X=1508798 $Y=1351110
X959 14450 13959 14675 14732 24 25 MXI2X1 $T=1508800 1473130 1 0 $X=1508798 $Y=1469190
X960 14255 13885 14694 14733 24 25 MXI2X1 $T=1508800 1532170 1 0 $X=1508798 $Y=1528230
X961 14467 13885 14700 14741 24 25 MXI2X1 $T=1509260 1539550 1 0 $X=1509258 $Y=1535610
X962 13850 497 14573 14668 24 25 MXI2X1 $T=1512480 1369810 1 180 $X=1509260 $Y=1369558
X963 14356 14131 14559 14649 24 25 MXI2X1 $T=1512480 1414090 1 180 $X=1509260 $Y=1413838
X964 14255 497 14691 14664 24 25 MXI2X1 $T=1512480 1502650 0 180 $X=1509260 $Y=1498710
X965 472 520 14730 14688 24 25 MXI2X1 $T=1509720 1362430 1 0 $X=1509718 $Y=1358490
X966 14467 13959 14771 14729 24 25 MXI2X1 $T=1509720 1517410 0 0 $X=1509718 $Y=1517158
X967 14421 14358 14738 14746 24 25 MXI2X1 $T=1511100 1428850 1 0 $X=1511098 $Y=1424910
X968 14255 14131 14773 14687 24 25 MXI2X1 $T=1517540 1480510 0 0 $X=1517538 $Y=1480258
X969 14255 14273 14699 14774 24 25 MXI2X1 $T=1517540 1502650 1 0 $X=1517538 $Y=1498710
X970 13850 14273 14695 14736 24 25 MXI2X1 $T=1520760 1369810 1 180 $X=1517540 $Y=1369558
X971 14356 13959 14766 14689 24 25 MXI2X1 $T=1520760 1414090 1 180 $X=1517540 $Y=1413838
X972 14421 14168 14682 14698 24 25 MXI2X1 $T=1520760 1443610 1 180 $X=1517540 $Y=1443358
X973 14467 14131 14758 14665 24 25 MXI2X1 $T=1519840 1502650 0 0 $X=1519838 $Y=1502398
X974 13850 14168 14783 14751 24 25 MXI2X1 $T=1523060 1391950 1 180 $X=1519840 $Y=1391698
X975 14450 14273 14784 14739 24 25 MXI2X1 $T=1523060 1473130 1 180 $X=1519840 $Y=1472878
X976 14230 14318 14785 14693 24 25 MXI2X1 $T=1523060 1510030 0 180 $X=1519840 $Y=1506090
X977 14421 13959 14789 14735 24 25 MXI2X1 $T=1521220 1450990 0 0 $X=1521218 $Y=1450738
X978 14467 14168 14953 14843 24 25 MXI2X1 $T=1523520 1502650 0 0 $X=1523518 $Y=1502398
X979 14255 14168 14850 14860 24 25 MXI2X1 $T=1523980 1502650 1 0 $X=1523978 $Y=1498710
X980 14467 14859 14841 14834 24 25 MXI2X1 $T=1527200 1487890 1 180 $X=1523980 $Y=1487638
X981 14450 14318 14750 14767 24 25 MXI2X1 $T=1527660 1465750 1 180 $X=1524440 $Y=1465498
X982 14421 14273 14737 14760 24 25 MXI2X1 $T=1524900 1414090 0 0 $X=1524898 $Y=1413838
X983 14450 14168 14845 14747 24 25 MXI2X1 $T=1528120 1443610 1 180 $X=1524900 $Y=1443358
X984 14421 14318 14761 14674 24 25 MXI2X1 $T=1528580 1436230 0 180 $X=1525360 $Y=1432290
X985 13850 14318 14867 14871 24 25 MXI2X1 $T=1526280 1384570 0 0 $X=1526278 $Y=1384318
X986 14450 14358 14772 14686 24 25 MXI2X1 $T=1529500 1473130 1 180 $X=1526280 $Y=1472878
X987 471 527 14855 14880 24 25 MXI2X1 $T=1526740 1355050 1 0 $X=1526738 $Y=1351110
X988 471 529 14742 14821 24 25 MXI2X1 $T=1526740 1362430 0 0 $X=1526738 $Y=1362178
X989 13850 14358 14927 14840 24 25 MXI2X1 $T=1526740 1384570 1 0 $X=1526738 $Y=1380630
X990 14356 14168 14933 14848 24 25 MXI2X1 $T=1526740 1399330 1 0 $X=1526738 $Y=1395390
X991 14356 14318 14864 14863 24 25 MXI2X1 $T=1526740 1406710 0 0 $X=1526738 $Y=1406458
X992 14854 335 14865 14925 24 25 MXI2X1 $T=1526740 1436230 0 0 $X=1526738 $Y=1435978
X993 14230 14859 14878 14836 24 25 MXI2X1 $T=1533180 1465750 1 180 $X=1529960 $Y=1465498
X994 14356 14358 14928 14842 24 25 MXI2X1 $T=1530880 1414090 0 0 $X=1530878 $Y=1413838
X995 14882 334 14916 14925 24 25 MXI2X1 $T=1531340 1443610 0 0 $X=1531338 $Y=1443358
X996 545 10382 14923 14937 24 25 MXI2X1 $T=1532260 1362430 1 0 $X=1532258 $Y=1358490
X997 14922 10297 14857 14941 24 25 MXI2X1 $T=1533180 1450990 0 0 $X=1533178 $Y=1450738
X998 14255 14358 14875 14976 24 25 MXI2X1 $T=1533180 1495270 0 0 $X=1533178 $Y=1495018
X999 546 10382 14943 14960 24 25 MXI2X1 $T=1534560 1377190 1 0 $X=1534558 $Y=1373250
X1000 14935 10297 14866 14957 24 25 MXI2X1 $T=1534560 1458370 1 0 $X=1534558 $Y=1454430
X1001 14467 14358 14926 14837 24 25 MXI2X1 $T=1535020 1517410 0 0 $X=1535018 $Y=1517158
X1002 14255 14859 14868 14930 24 25 MXI2X1 $T=1538240 1473130 1 180 $X=1535020 $Y=1472878
X1003 14450 14859 14939 14853 24 25 MXI2X1 $T=1539620 1414090 1 180 $X=1536400 $Y=1413838
X1004 472 529 15055 558 24 25 MXI2X1 $T=1541460 1355050 0 0 $X=1541458 $Y=1354798
X1005 14230 553 15058 15057 24 25 MXI2X1 $T=1541460 1480510 0 0 $X=1541458 $Y=1480258
X1006 14467 553 15034 15059 24 25 MXI2X1 $T=1541460 1487890 1 0 $X=1541458 $Y=1483950
X1007 546 562 15094 15067 24 25 MXI2X1 $T=1542840 1377190 1 0 $X=1542838 $Y=1373250
X1008 13891 553 15044 15064 24 25 MXI2X1 $T=1542840 1391950 0 0 $X=1542838 $Y=1391698
X1009 560 563 15029 15061 24 25 MXI2X1 $T=1542840 1414090 1 0 $X=1542838 $Y=1410150
X1010 560 562 14984 15062 24 25 MXI2X1 $T=1542840 1414090 0 0 $X=1542838 $Y=1413838
X1011 13836 553 15081 14973 24 25 MXI2X1 $T=1542840 1450990 1 0 $X=1542838 $Y=1447050
X1012 14922 563 15048 15091 24 25 MXI2X1 $T=1542840 1450990 0 0 $X=1542838 $Y=1450738
X1013 14450 553 15065 14952 24 25 MXI2X1 $T=1544220 1421470 0 0 $X=1544218 $Y=1421218
X1014 14356 14859 15071 15149 24 25 MXI2X1 $T=1548360 1399330 0 0 $X=1548358 $Y=1399078
X1015 14421 14859 15072 15139 24 25 MXI2X1 $T=1548360 1428850 0 0 $X=1548358 $Y=1428598
X1016 13836 14859 15135 15031 24 25 MXI2X1 $T=1548360 1436230 0 0 $X=1548358 $Y=1435978
X1017 15129 549 15032 14935 24 25 MXI2X1 $T=1551580 1458370 1 180 $X=1548360 $Y=1458118
X1018 15056 562 15131 15175 24 25 MXI2X1 $T=1552040 1406710 1 0 $X=1552038 $Y=1402770
X1019 13877 14859 15078 15045 24 25 MXI2X1 $T=1555260 1480510 0 180 $X=1552040 $Y=1476570
X1020 14032 14859 15053 15153 24 25 MXI2X1 $T=1558020 1487890 1 180 $X=1554800 $Y=1487638
X1021 577 562 15178 15235 24 25 MXI2X1 $T=1559400 1384570 0 0 $X=1559398 $Y=1384318
X1022 15056 563 15171 15238 24 25 MXI2X1 $T=1559400 1406710 0 0 $X=1559398 $Y=1406458
X1023 15187 563 15040 15245 24 25 MXI2X1 $T=1559400 1450990 0 0 $X=1559398 $Y=1450738
X1024 15187 562 15177 15236 24 25 MXI2X1 $T=1559400 1458370 0 0 $X=1559398 $Y=1458118
X1025 578 562 15173 15263 24 25 MXI2X1 $T=1560320 1465750 0 0 $X=1560318 $Y=1465498
X1026 15194 549 15233 15270 24 25 MXI2X1 $T=1560320 1495270 1 0 $X=1560318 $Y=1491330
X1027 15241 549 15163 577 24 25 MXI2X1 $T=1563540 1384570 0 180 $X=1560320 $Y=1380630
X1028 13850 14859 15239 15243 24 25 MXI2X1 $T=1560780 1377190 0 0 $X=1560778 $Y=1376938
X1029 13877 553 15257 15249 24 25 MXI2X1 $T=1561240 1465750 1 0 $X=1561238 $Y=1461810
X1030 13894 14859 15136 15228 24 25 MXI2X1 $T=1564460 1450990 0 180 $X=1561240 $Y=1447050
X1031 14421 553 15256 15267 24 25 MXI2X1 $T=1561700 1421470 1 0 $X=1561698 $Y=1417530
X1032 14032 553 15250 15231 24 25 MXI2X1 $T=1561700 1487890 1 0 $X=1561698 $Y=1483950
X1033 15247 549 14983 579 24 25 MXI2X1 $T=1564920 1399330 0 180 $X=1561700 $Y=1395390
X1034 583 563 14914 15260 24 25 MXI2X1 $T=1563080 1421470 0 0 $X=1563078 $Y=1421218
X1035 14255 553 15237 15253 24 25 MXI2X1 $T=1563540 1473130 0 0 $X=1563538 $Y=1472878
X1036 14356 553 15258 15320 24 25 MXI2X1 $T=1565840 1391950 1 0 $X=1565838 $Y=1388010
X1037 15268 575 15230 579 24 25 MXI2X1 $T=1569060 1399330 1 180 $X=1565840 $Y=1399078
X1038 15269 575 15261 15242 24 25 MXI2X1 $T=1569060 1436230 0 180 $X=1565840 $Y=1432290
X1039 13850 553 15264 15318 24 25 MXI2X1 $T=1566760 1384570 1 0 $X=1566758 $Y=1380630
X1040 13844 14859 15271 15176 24 25 MXI2X1 $T=1567680 1406710 0 0 $X=1567678 $Y=1406458
X1041 15281 549 15192 15242 24 25 MXI2X1 $T=1570900 1443610 0 180 $X=1567680 $Y=1439670
X1042 13894 553 15259 15324 24 25 MXI2X1 $T=1570440 1450990 1 0 $X=1570438 $Y=1447050
X1043 15322 549 15186 578 24 25 MXI2X1 $T=1573660 1465750 0 180 $X=1570440 $Y=1461810
X1044 13844 553 15328 15248 24 25 MXI2X1 $T=1572280 1406710 0 0 $X=1572278 $Y=1406458
X1045 583 562 15333 15332 24 25 MXI2X1 $T=1572280 1421470 0 0 $X=1572278 $Y=1421218
X1046 15270 562 15321 15337 24 25 MXI2X1 $T=1573200 1473130 1 0 $X=1573198 $Y=1469190
X1047 9745 25 35 24 9736 AND2X2 $T=1093420 1391950 1 0 $X=1093418 $Y=1388010
X1048 9927 25 9932 24 66 AND2X2 $T=1105380 1399330 1 0 $X=1105378 $Y=1395390
X1049 10031 25 10039 24 10065 AND2X2 $T=1115500 1406710 1 0 $X=1115498 $Y=1402770
X1050 10367 25 9939 24 10396 AND2X2 $T=1150920 1421470 0 0 $X=1150918 $Y=1421218
X1051 10466 25 10376 24 10494 AND2X2 $T=1151380 1355050 0 0 $X=1151378 $Y=1354798
X1052 119 25 141 24 10735 AND2X2 $T=1172080 1377190 0 0 $X=1172078 $Y=1376938
X1053 10931 25 69 24 10775 AND2X2 $T=1186800 1450990 0 0 $X=1186798 $Y=1450738
X1054 11299 25 10954 24 11387 AND2X2 $T=1216240 1399330 1 0 $X=1216238 $Y=1395390
X1055 11441 25 11454 24 11332 AND2X2 $T=1222220 1399330 0 180 $X=1220380 $Y=1395390
X1056 11301 25 189 24 11350 AND2X2 $T=1222680 1406710 0 180 $X=1220840 $Y=1402770
X1057 11508 25 11577 24 11644 AND2X2 $T=1231420 1369810 0 0 $X=1231418 $Y=1369558
X1058 124 25 10931 24 12030 AND2X2 $T=1259940 1524790 1 0 $X=1259938 $Y=1520850
X1059 111 25 10931 24 12027 AND2X2 $T=1259940 1532170 0 0 $X=1259938 $Y=1531918
X1060 12117 25 12077 24 12203 AND2X2 $T=1271900 1399330 0 0 $X=1271898 $Y=1399078
X1061 12030 25 12099 24 12118 AND2X2 $T=1271900 1524790 1 0 $X=1271898 $Y=1520850
X1062 12217 25 12210 24 12178 AND2X2 $T=1276040 1473130 0 180 $X=1274200 $Y=1469190
X1063 12230 25 12203 24 12346 AND2X2 $T=1279260 1399330 0 0 $X=1279258 $Y=1399078
X1064 12693 25 12685 24 329 AND2X2 $T=1315140 1362430 0 180 $X=1313300 $Y=1358490
X1065 12778 25 12685 24 333 AND2X2 $T=1322040 1362430 1 180 $X=1320200 $Y=1362178
X1066 12819 25 12685 24 341 AND2X2 $T=1326640 1362430 0 180 $X=1324800 $Y=1358490
X1067 12736 25 12676 24 12840 AND2X2 $T=1327560 1369810 1 0 $X=1327558 $Y=1365870
X1068 12894 25 12819 24 368 AND2X2 $T=1334000 1355050 0 0 $X=1333998 $Y=1354798
X1069 12894 25 12778 24 369 AND2X2 $T=1334460 1362430 1 0 $X=1334458 $Y=1358490
X1070 12894 25 12693 24 371 AND2X2 $T=1335840 1355050 0 0 $X=1335838 $Y=1354798
X1071 12670 25 12916 24 12894 AND2X2 $T=1339060 1362430 1 180 $X=1337220 $Y=1362178
X1072 12894 25 12793 24 355 AND2X2 $T=1337680 1355050 0 0 $X=1337678 $Y=1354798
X1073 12916 25 12676 24 12948 AND2X2 $T=1337680 1362430 1 0 $X=1337678 $Y=1358490
X1074 12884 25 12676 24 13015 AND2X2 $T=1340440 1369810 1 0 $X=1340438 $Y=1365870
X1075 12676 25 12901 24 13018 AND2X2 $T=1340900 1362430 1 0 $X=1340898 $Y=1358490
X1076 12670 25 12901 24 13040 AND2X2 $T=1344120 1362430 1 0 $X=1344118 $Y=1358490
X1077 12670 25 12884 24 13048 AND2X2 $T=1345960 1362430 0 0 $X=1345958 $Y=1362178
X1078 13040 25 12793 24 411 AND2X2 $T=1364820 1362430 1 0 $X=1364818 $Y=1358490
X1079 13040 25 12778 24 423 AND2X2 $T=1373560 1362430 1 0 $X=1373558 $Y=1358490
X1080 13040 25 12819 24 438 AND2X2 $T=1382760 1362430 1 0 $X=1382758 $Y=1358490
X1081 13040 25 12693 24 439 AND2X2 $T=1385980 1362430 1 0 $X=1385978 $Y=1358490
X1082 13048 25 12819 24 452 AND2X2 $T=1400700 1362430 1 0 $X=1400698 $Y=1358490
X1083 13048 25 12793 24 462 AND2X2 $T=1405760 1362430 1 0 $X=1405758 $Y=1358490
X1084 13048 25 12778 24 463 AND2X2 $T=1418640 1362430 1 180 $X=1416800 $Y=1362178
X1085 13048 25 12693 24 464 AND2X2 $T=1420480 1362430 0 0 $X=1420478 $Y=1362178
X1086 12840 25 12693 24 483 AND2X2 $T=1431060 1362430 1 0 $X=1431058 $Y=1358490
X1087 12840 25 12793 24 476 AND2X2 $T=1434740 1362430 1 0 $X=1434738 $Y=1358490
X1088 12840 25 12819 24 488 AND2X2 $T=1439340 1362430 1 0 $X=1439338 $Y=1358490
X1089 12840 25 12778 24 489 AND2X2 $T=1445320 1362430 1 0 $X=1445318 $Y=1358490
X1090 13015 25 12793 24 501 AND2X2 $T=1450840 1362430 1 0 $X=1450838 $Y=1358490
X1091 13015 25 12693 24 505 AND2X2 $T=1456360 1362430 1 0 $X=1456358 $Y=1358490
X1092 13015 25 12778 24 510 AND2X2 $T=1462340 1362430 1 0 $X=1462338 $Y=1358490
X1093 13015 25 12819 24 515 AND2X2 $T=1464640 1355050 1 0 $X=1464638 $Y=1351110
X1094 12948 25 12819 24 520 AND2X2 $T=1479360 1362430 1 0 $X=1479358 $Y=1358490
X1095 12948 25 12778 24 517 AND2X2 $T=1481660 1362430 1 0 $X=1481658 $Y=1358490
X1096 12948 25 12693 24 509 AND2X2 $T=1484420 1362430 1 0 $X=1484418 $Y=1358490
X1097 12948 25 12793 24 523 AND2X2 $T=1486720 1362430 1 0 $X=1486718 $Y=1358490
X1098 13018 25 12793 24 527 AND2X2 $T=1489480 1355050 0 0 $X=1489478 $Y=1354798
X1099 13018 25 12778 24 529 AND2X2 $T=1490860 1362430 1 0 $X=1490858 $Y=1358490
X1100 13018 25 12693 24 528 AND2X2 $T=1491780 1355050 0 0 $X=1491778 $Y=1354798
X1101 10245 25 14836 24 14870 AND2X2 $T=1525820 1450990 0 0 $X=1525818 $Y=1450738
X1102 14821 25 14851 24 14950 AND2X2 $T=1531340 1369810 0 0 $X=1531338 $Y=1369558
X1103 10378 25 14853 24 14987 AND2X2 $T=1535940 1406710 0 0 $X=1535938 $Y=1406458
X1104 15041 25 15045 24 15073 AND2X2 $T=1544220 1480510 1 0 $X=1544218 $Y=1476570
X1105 10245 25 15060 24 15095 AND2X2 $T=1548820 1384570 1 0 $X=1548818 $Y=1380630
X1106 10245 25 15176 24 15130 AND2X2 $T=1557100 1406710 1 180 $X=1555260 $Y=1406458
X1107 15139 25 15142 24 15232 AND2X2 $T=1555720 1428850 0 0 $X=1555718 $Y=1428598
X1108 15153 25 15183 24 15184 AND2X2 $T=1558940 1480510 1 0 $X=1558938 $Y=1476570
X1109 15228 25 15191 24 15265 AND2X2 $T=1563080 1443610 1 0 $X=1563078 $Y=1439670
X1110 383 25 15320 24 15268 AND2X2 $T=1572740 1399330 0 0 $X=1572738 $Y=1399078
X1111 10737 10731 24 25 10724 AND2XL $T=1173920 1421470 1 180 $X=1172080 $Y=1421218
X1112 10762 10724 24 25 10779 AND2XL $T=1175760 1414090 1 0 $X=1175758 $Y=1410150
X1113 10742 10732 24 25 10848 AND2XL $T=1178060 1399330 1 0 $X=1178058 $Y=1395390
X1114 10798 10779 24 25 10732 AND2XL $T=1181280 1399330 1 180 $X=1179440 $Y=1399078
X1115 158 10909 24 25 10731 AND2XL $T=1184960 1428850 0 180 $X=1183120 $Y=1424910
X1116 56 10931 24 25 10936 AND2XL $T=1185420 1458370 1 0 $X=1185418 $Y=1454430
X1117 10887 11042 24 25 10909 AND2XL $T=1194620 1436230 0 180 $X=1192780 $Y=1432290
X1118 78 10931 24 25 11084 AND2XL $T=1196000 1480510 1 0 $X=1195998 $Y=1476570
X1119 71 10931 24 25 11177 AND2XL $T=1198300 1495270 1 0 $X=1198298 $Y=1491330
X1120 11203 11110 24 25 11042 AND2XL $T=1200140 1443610 1 180 $X=1198300 $Y=1443358
X1121 143 10931 24 25 11129 AND2XL $T=1198760 1524790 1 0 $X=1198758 $Y=1520850
X1122 64 10931 24 25 11176 AND2XL $T=1199220 1480510 1 0 $X=1199218 $Y=1476570
X1123 67 10931 24 25 11068 AND2XL $T=1201980 1458370 1 180 $X=1200140 $Y=1458118
X1124 11211 11014 24 25 11086 AND2XL $T=1203820 1377190 1 180 $X=1201980 $Y=1376938
X1125 11178 10848 24 25 11301 AND2XL $T=1207040 1399330 1 0 $X=1207038 $Y=1395390
X1126 117 10931 24 25 11128 AND2XL $T=1207040 1510030 0 0 $X=1207038 $Y=1509778
X1127 11227 11246 24 25 11110 AND2XL $T=1210720 1458370 1 180 $X=1208880 $Y=1458118
X1128 11317 11319 24 25 11309 AND2XL $T=1214860 1517410 0 180 $X=1213020 $Y=1513470
X1129 11316 11309 24 25 11367 AND2XL $T=1213940 1495270 0 0 $X=1213938 $Y=1495018
X1130 11383 11351 24 25 11246 AND2XL $T=1217160 1473130 1 180 $X=1215320 $Y=1472878
X1131 11362 11367 24 25 11351 AND2XL $T=1217160 1480510 0 0 $X=1217158 $Y=1480258
X1132 11313 11301 24 25 11485 AND2XL $T=1222220 1414090 1 0 $X=1222218 $Y=1410150
X1133 122 10931 24 25 11531 AND2XL $T=1232800 1524790 1 180 $X=1230960 $Y=1524538
X1134 11614 11601 24 25 11319 AND2XL $T=1234640 1510030 1 180 $X=1232800 $Y=1509778
X1135 108 10931 24 25 11627 AND2XL $T=1234640 1532170 1 0 $X=1234638 $Y=1528230
X1136 11647 11660 24 25 11683 AND2XL $T=1237400 1406710 0 0 $X=1237398 $Y=1406458
X1137 11073 11647 24 25 11509 AND2XL $T=1237400 1428850 1 0 $X=1237398 $Y=1424910
X1138 100 10931 24 25 11642 AND2XL $T=1241540 1532170 0 180 $X=1239700 $Y=1528230
X1139 11690 11666 24 25 11601 AND2XL $T=1243380 1510030 1 180 $X=1241540 $Y=1509778
X1140 11775 11683 24 25 11892 AND2XL $T=1247520 1399330 0 0 $X=1247518 $Y=1399078
X1141 88 10931 24 25 11809 AND2XL $T=1247520 1532170 1 0 $X=1247518 $Y=1528230
X1142 11739 11760 24 25 11666 AND2XL $T=1250280 1510030 0 180 $X=1248440 $Y=1506090
X1143 11918 11891 24 25 11760 AND2XL $T=1251660 1510030 1 180 $X=1249820 $Y=1509778
X1144 95 10931 24 25 11919 AND2XL $T=1255800 1532170 1 180 $X=1253960 $Y=1531918
X1145 12014 11944 24 25 11891 AND2XL $T=1257640 1517410 0 180 $X=1255800 $Y=1513470
X1146 11925 11892 24 25 12019 AND2XL $T=1257180 1399330 0 0 $X=1257178 $Y=1399078
X1147 65 10931 24 25 12038 AND2XL $T=1260860 1524790 0 0 $X=1260858 $Y=1524538
X1148 12053 12019 24 25 12077 AND2XL $T=1264080 1399330 0 0 $X=1264078 $Y=1399078
X1149 12173 12105 24 25 11944 AND2XL $T=1269600 1510030 1 180 $X=1267760 $Y=1509778
X1150 12228 12229 24 25 12105 AND2XL $T=1278340 1510030 1 180 $X=1276500 $Y=1509778
X1151 391 15324 24 25 15269 AND2XL $T=1574120 1436230 1 180 $X=1572280 $Y=1435978
X1152 10126 24 10013 10164 25 NAND2X1 $T=1128380 1436230 0 180 $X=1127000 $Y=1432290
X1153 10251 24 10234 10230 25 NAND2X1 $T=1132980 1473130 0 180 $X=1131600 $Y=1469190
X1154 10389 24 10455 10234 25 NAND2X1 $T=1150920 1473130 0 180 $X=1149540 $Y=1469190
X1155 142 24 144 10805 25 NAND2X1 $T=1172540 1355050 1 0 $X=1172538 $Y=1351110
X1156 141 24 119 10781 25 NAND2X1 $T=1174840 1458370 1 0 $X=1174838 $Y=1454430
X1157 150 24 10800 10872 25 NAND2X1 $T=1179900 1377190 0 0 $X=1179898 $Y=1376938
X1158 10875 24 10879 10917 25 NAND2X1 $T=1181740 1369810 0 0 $X=1181738 $Y=1369558
X1159 10925 24 155 10935 25 NAND2X1 $T=1185880 1362430 1 0 $X=1185878 $Y=1358490
X1160 10954 24 159 10815 25 NAND2X1 $T=1189560 1384570 0 180 $X=1188180 $Y=1380630
X1161 10954 24 11034 10893 25 NAND2X1 $T=1193700 1384570 0 180 $X=1192320 $Y=1380630
X1162 10971 24 10930 11058 25 NAND2X1 $T=1192780 1369810 0 0 $X=1192778 $Y=1369558
X1163 10954 24 167 11009 25 NAND2X1 $T=1194160 1384570 1 180 $X=1192780 $Y=1384318
X1164 11105 24 10970 10881 25 NAND2X1 $T=1197840 1487890 0 180 $X=1196460 $Y=1483950
X1165 10872 24 11016 11097 25 NAND2X1 $T=1196920 1377190 0 0 $X=1196918 $Y=1376938
X1166 11058 24 11078 11096 25 NAND2X1 $T=1197380 1369810 1 0 $X=1197378 $Y=1365870
X1167 10954 24 11074 11050 25 NAND2X1 $T=1198760 1384570 1 180 $X=1197380 $Y=1384318
X1168 11088 24 11107 11169 25 NAND2X1 $T=1198760 1362430 1 0 $X=1198758 $Y=1358490
X1169 178 24 10668 11088 25 NAND2X1 $T=1202440 1355050 0 180 $X=1201060 $Y=1351110
X1170 10954 24 11124 11212 25 NAND2X1 $T=1202900 1391950 1 0 $X=1202898 $Y=1388010
X1171 10954 24 177 11125 25 NAND2X1 $T=1204280 1384570 0 180 $X=1202900 $Y=1380630
X1172 10954 24 11182 11127 25 NAND2X1 $T=1204280 1384570 1 180 $X=1202900 $Y=1384318
X1173 11014 24 11236 11304 25 NAND2X1 $T=1208420 1384570 1 0 $X=1208418 $Y=1380630
X1174 10954 24 11221 11087 25 NAND2X1 $T=1209800 1384570 1 180 $X=1208420 $Y=1384318
X1175 11196 24 11254 11123 25 NAND2X1 $T=1209340 1502650 1 0 $X=1209338 $Y=1498710
X1176 11302 24 11262 11254 25 NAND2X1 $T=1211180 1502650 1 180 $X=1209800 $Y=1502398
X1177 10954 24 192 11343 25 NAND2X1 $T=1213020 1399330 1 0 $X=1213018 $Y=1395390
X1178 191 24 10767 11337 25 NAND2X1 $T=1213480 1384570 1 0 $X=1213478 $Y=1380630
X1179 11496 24 10751 11320 25 NAND2X1 $T=1215320 1391950 1 180 $X=1213940 $Y=1391698
X1180 198 24 11374 11445 25 NAND2X1 $T=1218540 1355050 1 0 $X=1218538 $Y=1351110
X1181 11337 24 11388 11448 25 NAND2X1 $T=1219460 1377190 0 0 $X=1219458 $Y=1376938
X1182 176 24 10797 11328 25 NAND2X1 $T=1222220 1369810 1 180 $X=1220840 $Y=1369558
X1183 11376 24 11452 11455 25 NAND2X1 $T=1223140 1428850 0 0 $X=1223138 $Y=1428598
X1184 10954 24 11453 11347 25 NAND2X1 $T=1224520 1436230 1 180 $X=1223140 $Y=1435978
X1185 196 24 11478 11370 25 NAND2X1 $T=1226360 1355050 1 180 $X=1224980 $Y=1354798
X1186 11513 24 11482 11472 25 NAND2X1 $T=1227740 1406710 0 180 $X=1226360 $Y=1402770
X1187 11522 24 11521 11537 25 NAND2X1 $T=1229580 1384570 0 0 $X=1229578 $Y=1384318
X1188 11498 24 10644 11577 25 NAND2X1 $T=1230500 1369810 1 0 $X=1230498 $Y=1365870
X1189 11534 24 11544 11582 25 NAND2X1 $T=1230960 1443610 1 0 $X=1230958 $Y=1439670
X1190 11580 24 11545 11380 25 NAND2X1 $T=1232340 1450990 1 180 $X=1230960 $Y=1450738
X1191 11580 24 11584 11344 25 NAND2X1 $T=1232800 1450990 0 180 $X=1231420 $Y=1447050
X1192 11530 24 10849 11649 25 NAND2X1 $T=1231880 1436230 1 0 $X=1231878 $Y=1432290
X1193 11580 24 11589 11444 25 NAND2X1 $T=1233260 1465750 1 180 $X=1231880 $Y=1465498
X1194 11620 24 10768 11602 25 NAND2X1 $T=1234640 1465750 0 180 $X=1233260 $Y=1461810
X1195 11580 24 11612 11619 25 NAND2X1 $T=1233720 1480510 1 0 $X=1233718 $Y=1476570
X1196 11534 24 11579 11657 25 NAND2X1 $T=1234180 1443610 0 0 $X=1234178 $Y=1443358
X1197 11587 24 11623 11663 25 NAND2X1 $T=1234640 1406710 1 0 $X=1234638 $Y=1402770
X1198 11593 24 11618 11639 25 NAND2X1 $T=1234640 1473130 1 0 $X=1234638 $Y=1469190
X1199 11580 24 11625 11488 25 NAND2X1 $T=1236020 1450990 1 180 $X=1234640 $Y=1450738
X1200 11650 24 11579 11544 25 NAND2X1 $T=1236940 1443610 0 180 $X=1235560 $Y=1439670
X1201 11580 24 11654 11392 25 NAND2X1 $T=1238320 1450990 0 180 $X=1236940 $Y=1447050
X1202 11580 24 11655 11609 25 NAND2X1 $T=1238320 1480510 0 180 $X=1236940 $Y=1476570
X1203 11652 24 11651 11682 25 NAND2X1 $T=1237400 1362430 1 0 $X=1237398 $Y=1358490
X1204 11662 24 10736 11653 25 NAND2X1 $T=1238780 1369810 1 180 $X=1237400 $Y=1369558
X1205 11659 24 11663 11670 25 NAND2X1 $T=1238320 1406710 1 0 $X=1238318 $Y=1402770
X1206 11320 24 11533 11734 25 NAND2X1 $T=1239240 1391950 0 0 $X=1239238 $Y=1391698
X1207 11652 24 11697 11787 25 NAND2X1 $T=1241540 1362430 0 0 $X=1241538 $Y=1362178
X1208 11768 24 11595 11656 25 NAND2X1 $T=1242920 1384570 0 180 $X=1241540 $Y=1380630
X1209 11602 24 11743 11795 25 NAND2X1 $T=1242920 1465750 0 0 $X=1242918 $Y=1465498
X1210 11744 24 10850 11805 25 NAND2X1 $T=1243380 1480510 0 0 $X=1243378 $Y=1480258
X1211 11793 24 11774 11868 25 NAND2X1 $T=1247060 1399330 1 0 $X=1247058 $Y=1395390
X1212 11689 24 11808 11799 25 NAND2X1 $T=1247980 1473130 1 0 $X=1247978 $Y=1469190
X1213 11580 24 11883 11747 25 NAND2X1 $T=1251200 1450990 1 180 $X=1249820 $Y=1450738
X1214 11580 24 11889 11900 25 NAND2X1 $T=1250740 1450990 1 0 $X=1250738 $Y=1447050
X1215 11805 24 11928 11962 25 NAND2X1 $T=1254420 1480510 1 0 $X=1254418 $Y=1476570
X1216 11948 24 10863 11937 25 NAND2X1 $T=1257180 1473130 0 0 $X=1257178 $Y=1472878
X1217 11580 24 12022 11936 25 NAND2X1 $T=1261780 1480510 0 180 $X=1260400 $Y=1476570
X1218 11937 24 11933 11884 25 NAND2X1 $T=1260860 1465750 1 0 $X=1260858 $Y=1461810
X1219 12048 24 11961 11913 25 NAND2X1 $T=1262700 1399330 1 180 $X=1261320 $Y=1399078
X1220 11580 24 12068 12094 25 NAND2X1 $T=1265460 1465750 1 0 $X=1265458 $Y=1461810
X1221 11580 24 12069 12087 25 NAND2X1 $T=1266380 1473130 0 0 $X=1266378 $Y=1472878
X1222 12073 24 12079 12088 25 NAND2X1 $T=1266380 1480510 0 0 $X=1266378 $Y=1480258
X1223 12059 24 12083 12116 25 NAND2X1 $T=1268680 1391950 1 0 $X=1268678 $Y=1388010
X1224 11580 24 12169 12096 25 NAND2X1 $T=1271440 1465750 0 180 $X=1270060 $Y=1461810
X1225 12201 24 10743 12184 25 NAND2X1 $T=1274660 1458370 0 0 $X=1274658 $Y=1458118
X1226 12222 24 11804 12176 25 NAND2X1 $T=1277880 1480510 0 0 $X=1277878 $Y=1480258
X1227 12315 24 11093 12235 25 NAND2X1 $T=1279720 1465750 1 180 $X=1278340 $Y=1465498
X1228 12235 24 12262 12250 25 NAND2X1 $T=1278800 1458370 0 0 $X=1278798 $Y=1458118
X1229 12176 24 12242 12199 25 NAND2X1 $T=1278800 1473130 1 0 $X=1278798 $Y=1469190
X1230 101 24 12366 12628 25 NAND2X1 $T=1307320 1450990 0 0 $X=1307318 $Y=1450738
X1231 12736 24 12670 12673 25 NAND2X1 $T=1317900 1362430 1 180 $X=1316520 $Y=1362178
X1232 14865 24 14844 14072 25 NAND2X1 $T=1526280 1443610 0 180 $X=1524900 $Y=1439670
X1233 14866 24 14856 14418 25 NAND2X1 $T=1528580 1458370 0 180 $X=1527200 $Y=1454430
X1234 14938 24 14857 14589 25 NAND2X1 $T=1528580 1465750 0 180 $X=1527200 $Y=1461810
X1235 14914 24 14881 14681 25 NAND2X1 $T=1531800 1428850 0 180 $X=1530420 $Y=1424910
X1236 14916 24 14931 14075 25 NAND2X1 $T=1534100 1443610 1 0 $X=1534098 $Y=1439670
X1237 14943 24 14946 14073 25 NAND2X1 $T=1537320 1377190 1 180 $X=1535940 $Y=1376938
X1238 14984 24 14944 14588 25 NAND2X1 $T=1537320 1428850 1 180 $X=1535940 $Y=1428598
X1239 14923 24 14954 14183 25 NAND2X1 $T=1536400 1362430 0 0 $X=1536398 $Y=1362178
X1240 14983 24 14951 14625 25 NAND2X1 $T=1537780 1399330 0 180 $X=1536400 $Y=1395390
X1241 15029 24 14972 14524 25 NAND2X1 $T=1540080 1414090 0 180 $X=1538700 $Y=1410150
X1242 15032 24 14970 14417 25 NAND2X1 $T=1540080 1465750 1 180 $X=1538700 $Y=1465498
X1243 557 24 14985 14354 25 NAND2X1 $T=1542380 1369810 0 180 $X=1541000 $Y=1365870
X1244 15040 24 15033 14067 25 NAND2X1 $T=1543760 1465750 0 180 $X=1542380 $Y=1461810
X1245 15131 24 15047 14117 25 NAND2X1 $T=1545600 1406710 0 180 $X=1544220 $Y=1402770
X1246 15048 24 15054 14516 25 NAND2X1 $T=1544680 1502650 0 0 $X=1544678 $Y=1502398
X1247 15094 24 15126 14074 25 NAND2X1 $T=1550200 1377190 1 0 $X=1550198 $Y=1373250
X1248 15173 24 15143 14577 25 NAND2X1 $T=1554800 1473130 1 180 $X=1553420 $Y=1472878
X1249 15233 24 15144 14165 25 NAND2X1 $T=1554800 1502650 1 180 $X=1553420 $Y=1502398
X1250 572 24 15156 14648 25 NAND2X1 $T=1556180 1362430 1 180 $X=1554800 $Y=1362178
X1251 15163 24 15157 14643 25 NAND2X1 $T=1556180 1384570 0 180 $X=1554800 $Y=1380630
X1252 15186 24 15093 14521 25 NAND2X1 $T=1556180 1465750 1 180 $X=1554800 $Y=1465498
X1253 15171 24 15160 14146 25 NAND2X1 $T=1556640 1414090 0 180 $X=1555260 $Y=1410150
X1254 15192 24 15150 13876 25 NAND2X1 $T=1556640 1450990 0 180 $X=1555260 $Y=1447050
X1255 15177 24 15162 14065 25 NAND2X1 $T=1556640 1458370 1 180 $X=1555260 $Y=1458118
X1256 15178 24 15172 14582 25 NAND2X1 $T=1559400 1384570 1 180 $X=1558020 $Y=1384318
X1257 15230 24 15193 14576 25 NAND2X1 $T=1561700 1399330 1 180 $X=1560320 $Y=1399078
X1258 15261 24 15227 14185 25 NAND2X1 $T=1562160 1436230 1 180 $X=1560780 $Y=1435978
X1259 15321 24 15190 14127 25 NAND2X1 $T=1570440 1473130 1 180 $X=1569060 $Y=1472878
X1260 15333 24 15285 14626 25 NAND2X1 $T=1572740 1428850 1 180 $X=1571360 $Y=1428598
X1261 12370 12474 12468 11960 12404 12342 11470 24 25 12331 SDFFNSRXL $T=1294440 1532170 0 180 $X=1282480 $Y=1528230
X1262 12370 12382 12389 11960 12404 12342 12474 24 25 12520 SDFFNSRXL $T=1286160 1524790 0 0 $X=1286158 $Y=1524538
X1263 12370 12388 12395 11960 296 12497 12513 24 25 12516 SDFFNSRXL $T=1286620 1539550 1 0 $X=1286618 $Y=1535610
X1264 289 12348 12378 229 10062 12506 12336 24 25 319 SDFFNSRXL $T=1287080 1369810 1 0 $X=1287078 $Y=1365870
X1265 289 12391 12397 229 10062 12507 12365 24 25 12521 SDFFNSRXL $T=1287080 1384570 1 0 $X=1287078 $Y=1380630
X1266 11874 12392 12377 12113 12404 12508 12479 24 25 12594 SDFFNSRXL $T=1287080 1450990 1 0 $X=1287078 $Y=1447050
X1267 12478 12413 12501 12113 12404 12398 12369 24 25 12383 SDFFNSRXL $T=1299040 1421470 1 180 $X=1287080 $Y=1421218
X1268 11874 12479 12502 12113 12404 12399 11922 24 25 12385 SDFFNSRXL $T=1299040 1465750 0 180 $X=1287080 $Y=1461810
X1269 12478 12365 12527 229 12404 12462 12413 24 25 12410 SDFFNSRXL $T=1301800 1406710 0 180 $X=1289840 $Y=1402770
X1270 11874 290 12464 12113 12404 12560 12496 24 25 12569 SDFFNSRXL $T=1290300 1458370 0 0 $X=1290298 $Y=1458118
X1271 12054 12496 12503 12113 12404 12615 12486 24 25 12626 SDFFNSRXL $T=1295820 1480510 0 0 $X=1295818 $Y=1480258
X1272 12370 12526 12561 11960 296 12497 12388 24 25 12669 SDFFNSRXL $T=1299040 1539550 1 0 $X=1299038 $Y=1535610
X1273 12478 12562 12563 229 296 12462 12601 24 25 12680 SDFFNSRXL $T=1299960 1406710 0 0 $X=1299958 $Y=1406458
X1274 12370 12567 12575 11960 321 12342 12618 24 25 12677 SDFFNSRXL $T=1300880 1524790 0 0 $X=1300878 $Y=1524538
X1275 11874 12573 12522 12113 322 12508 12515 24 25 12710 SDFFNSRXL $T=1301340 1443610 0 0 $X=1301338 $Y=1443358
X1276 11874 12574 12579 12113 12404 12560 12227 24 25 12697 SDFFNSRXL $T=1301340 1458370 1 0 $X=1301338 $Y=1454430
X1277 11874 12582 12589 12113 296 12399 12583 24 25 12689 SDFFNSRXL $T=1302260 1465750 1 0 $X=1302258 $Y=1461810
X1278 12054 12591 12598 12113 322 12678 12403 24 25 12690 SDFFNSRXL $T=1302720 1487890 1 0 $X=1302718 $Y=1483950
X1279 12411 12486 12523 12113 12404 12679 12564 24 25 12728 SDFFNSRXL $T=1302720 1487890 0 0 $X=1302718 $Y=1487638
X1280 289 12578 12607 229 325 12683 12391 24 25 12719 SDFFNSRXL $T=1303640 1377190 0 0 $X=1303638 $Y=1376938
X1281 12411 12599 12605 11960 321 12684 12637 24 25 12791 SDFFNSRXL $T=1303640 1502650 0 0 $X=1303638 $Y=1502398
X1282 12478 12672 12674 229 12641 12462 12562 24 25 12577 SDFFNSRXL $T=1315600 1406710 0 180 $X=1303640 $Y=1402770
X1283 289 320 12585 229 324 12683 12166 24 25 12714 SDFFNSRXL $T=1304100 1384570 1 0 $X=1304098 $Y=1380630
X1284 12478 12601 12609 12113 321 12687 12602 24 25 12706 SDFFNSRXL $T=1304100 1421470 1 0 $X=1304098 $Y=1417530
X1285 12478 12581 12588 12113 12404 12688 12573 24 25 12727 SDFFNSRXL $T=1304100 1436230 0 0 $X=1304098 $Y=1435978
X1286 12054 12604 12612 11960 322 12684 11806 24 25 12695 SDFFNSRXL $T=1304100 1495270 0 0 $X=1304098 $Y=1495018
X1287 12411 12564 12592 11960 12404 12684 12488 24 25 12784 SDFFNSRXL $T=1304100 1502650 1 0 $X=1304098 $Y=1498710
X1288 12370 12611 12596 11960 322 12692 12593 24 25 12703 SDFFNSRXL $T=1304560 1546930 0 0 $X=1304558 $Y=1546678
X1289 11874 12515 12620 12113 327 12508 12702 24 25 12731 SDFFNSRXL $T=1305020 1450990 1 0 $X=1305018 $Y=1447050
X1290 12054 12629 12631 12113 327 12615 12591 24 25 12712 SDFFNSRXL $T=1307780 1480510 0 0 $X=1307778 $Y=1480258
X1291 12370 12488 12632 11960 12404 12721 12382 24 25 12732 SDFFNSRXL $T=1307780 1524790 1 0 $X=1307778 $Y=1520850
X1292 12370 12513 12576 11960 321 12342 12606 24 25 12786 SDFFNSRXL $T=1307780 1532170 0 0 $X=1307778 $Y=1531918
X1293 12054 12630 12638 12113 296 12615 12629 24 25 12711 SDFFNSRXL $T=1308240 1473130 0 0 $X=1308238 $Y=1472878
X1294 12370 12633 12639 11960 296 12497 12611 24 25 12730 SDFFNSRXL $T=1308240 1546930 1 0 $X=1308238 $Y=1542990
X1295 12411 12637 12640 11960 322 12684 12642 24 25 12742 SDFFNSRXL $T=1308700 1510030 0 0 $X=1308698 $Y=1509778
X1296 12478 12737 12571 12113 322 12398 12603 24 25 12634 SDFFNSRXL $T=1321120 1421470 1 180 $X=1309160 $Y=1421218
X1297 12370 12686 12691 11960 296 12721 12715 24 25 12808 SDFFNSRXL $T=1313300 1517410 0 0 $X=1313298 $Y=1517158
X1298 289 12696 12700 229 327 12507 12774 24 25 12821 SDFFNSRXL $T=1314680 1384570 0 0 $X=1314678 $Y=1384318
X1299 289 12699 12705 229 321 12506 12696 24 25 12824 SDFFNSRXL $T=1315140 1377190 1 0 $X=1315138 $Y=1373250
X1300 12370 12642 12713 11960 322 12721 12633 24 25 12708 SDFFNSRXL $T=1315600 1517410 1 0 $X=1315598 $Y=1513470
X1301 318 332 12716 229 321 12818 331 24 25 350 SDFFNSRXL $T=1316060 1355050 1 0 $X=1316058 $Y=1351110
X1302 12370 12715 12722 11960 337 12805 12738 24 25 12833 SDFFNSRXL $T=1316520 1561690 1 0 $X=1316518 $Y=1557750
X1303 289 12835 12744 229 327 12683 12699 24 25 12723 SDFFNSRXL $T=1330320 1377190 1 180 $X=1318360 $Y=1376938
X1304 12411 12781 12789 11960 337 12684 12686 24 25 12878 SDFFNSRXL $T=1320660 1510030 0 0 $X=1320658 $Y=1509778
X1305 12478 12830 12826 12113 321 12787 12777 24 25 12745 SDFFNSRXL $T=1332620 1443610 0 180 $X=1320660 $Y=1439670
X1306 12597 12872 12746 12113 322 12560 12617 24 25 12772 SDFFNSRXL $T=1333080 1458370 0 180 $X=1321120 $Y=1454430
X1307 289 12774 12785 229 321 12507 12780 24 25 12834 SDFFNSRXL $T=1321580 1391950 0 0 $X=1321578 $Y=1391698
X1308 12478 338 12775 12113 322 12687 12737 24 25 12838 SDFFNSRXL $T=1321580 1414090 0 0 $X=1321578 $Y=1413838
X1309 12597 12776 12794 12113 337 12615 12630 24 25 12885 SDFFNSRXL $T=1321580 1473130 0 0 $X=1321578 $Y=1472878
X1310 12597 12877 12743 12113 321 12615 12776 24 25 12783 SDFFNSRXL $T=1333540 1480510 0 180 $X=1321580 $Y=1476570
X1311 12478 12777 12800 12113 12404 12688 12796 24 25 12889 SDFFNSRXL $T=1322040 1436230 1 0 $X=1322038 $Y=1432290
X1312 12478 12796 12803 12113 12641 12398 12627 24 25 12908 SDFFNSRXL $T=1322500 1428850 1 0 $X=1322498 $Y=1424910
X1313 12370 12799 12804 11960 348 12342 12801 24 25 13034 SDFFNSRXL $T=1322500 1532170 0 0 $X=1322498 $Y=1531918
X1314 12957 12738 12881 11960 337 12805 12795 24 25 12792 SDFFNSRXL $T=1334460 1554310 1 180 $X=1322500 $Y=1554058
X1315 12597 12898 12843 11960 321 12679 12604 24 25 12741 SDFFNSRXL $T=1335840 1495270 0 180 $X=1323880 $Y=1491330
X1316 12411 12896 12909 11960 348 12721 12781 24 25 12815 SDFFNSRXL $T=1337220 1517410 1 180 $X=1325260 $Y=1517158
X1317 12597 12827 12831 12113 348 12925 12877 24 25 12964 SDFFNSRXL $T=1326640 1473130 1 0 $X=1326638 $Y=1469190
X1318 12597 12842 12844 12113 348 12678 12886 24 25 12973 SDFFNSRXL $T=1329400 1487890 0 0 $X=1329398 $Y=1487638
X1319 12411 12873 12879 11960 348 12974 12799 24 25 13017 SDFFNSRXL $T=1330780 1546930 1 0 $X=1330778 $Y=1542990
X1320 12597 12883 12888 11960 348 12684 12904 24 25 13022 SDFFNSRXL $T=1332160 1502650 0 0 $X=1332158 $Y=1502398
X1321 12597 12886 12895 11960 12641 12679 12883 24 25 13024 SDFFNSRXL $T=1332620 1495270 0 0 $X=1332618 $Y=1495018
X1322 12597 12590 12911 12113 12641 12615 12842 24 25 12950 SDFFNSRXL $T=1334460 1480510 0 0 $X=1334458 $Y=1480258
X1323 12411 12904 12914 11960 375 13025 12937 24 25 13036 SDFFNSRXL $T=1334460 1510030 0 0 $X=1334458 $Y=1509778
X1324 12478 13027 12841 12113 337 12688 12830 24 25 12902 SDFFNSRXL $T=1346420 1436230 0 180 $X=1334460 $Y=1432290
X1325 366 12782 12920 229 378 12507 12953 24 25 13049 SDFFNSRXL $T=1335380 1384570 0 0 $X=1335378 $Y=1384318
X1326 12478 12917 12921 229 348 12926 12836 24 25 13046 SDFFNSRXL $T=1335380 1399330 0 0 $X=1335378 $Y=1399078
X1327 12942 12924 12931 229 337 12926 12917 24 25 12912 SDFFNSRXL $T=1347800 1399330 0 180 $X=1335840 $Y=1395390
X1328 12597 12951 12906 12113 12641 12399 12907 24 25 12913 SDFFNSRXL $T=1347800 1465750 0 180 $X=1335840 $Y=1461810
X1329 12411 12937 12941 11960 12641 13042 12961 24 25 13050 SDFFNSRXL $T=1337220 1524790 0 0 $X=1337218 $Y=1524538
X1330 289 12947 12910 379 378 12506 12924 24 25 13094 SDFFNSRXL $T=1338140 1369810 0 0 $X=1338138 $Y=1369558
X1331 289 13030 13039 229 375 12683 12835 24 25 12939 SDFFNSRXL $T=1350100 1377190 1 180 $X=1338140 $Y=1376938
X1332 12942 12954 12963 12113 12641 12687 13035 24 25 13120 SDFFNSRXL $T=1338600 1414090 0 0 $X=1338598 $Y=1413838
X1333 12597 12927 12936 12113 12641 12560 12930 24 25 13103 SDFFNSRXL $T=1338600 1458370 0 0 $X=1338598 $Y=1458118
X1334 12942 12928 13045 12113 12641 12787 12949 24 25 12943 SDFFNSRXL $T=1350560 1443610 0 180 $X=1338600 $Y=1439670
X1335 12597 13055 12972 12113 375 12615 12951 24 25 12944 SDFFNSRXL $T=1350560 1480510 0 180 $X=1338600 $Y=1476570
X1336 12957 12945 13029 11960 375 12805 12956 24 25 12946 SDFFNSRXL $T=1350560 1561690 1 180 $X=1338600 $Y=1561438
X1337 12411 12961 12967 11960 348 13062 13061 24 25 13037 SDFFNSRXL $T=1339060 1539550 1 0 $X=1339058 $Y=1535610
X1338 289 377 12968 379 348 12818 13064 24 25 388 SDFFNSRXL $T=1339520 1355050 0 0 $X=1339518 $Y=1354798
X1339 12957 13014 12940 11960 12641 12692 12945 24 25 13110 SDFFNSRXL $T=1340900 1554310 1 0 $X=1340898 $Y=1550370
X1340 12597 13013 13041 12113 381 12678 12898 24 25 12975 SDFFNSRXL $T=1353320 1487890 1 180 $X=1341360 $Y=1487638
X1341 12942 12829 13020 229 12641 12462 12954 24 25 13105 SDFFNSRXL $T=1341820 1406710 0 0 $X=1341818 $Y=1406458
X1342 289 13117 12965 379 348 12506 12947 24 25 13016 SDFFNSRXL $T=1354700 1369810 0 180 $X=1342740 $Y=1365870
X1343 12597 362 13019 12113 12641 12678 13013 24 25 13132 SDFFNSRXL $T=1344120 1487890 1 0 $X=1344118 $Y=1483950
X1344 366 13137 13067 13102 348 12683 13030 24 25 13028 SDFFNSRXL $T=1357000 1384570 0 180 $X=1345040 $Y=1380630
X1345 12942 13035 13093 13102 375 12398 13108 24 25 13140 SDFFNSRXL $T=1349640 1421470 0 0 $X=1349638 $Y=1421218
X1346 12411 13186 13167 11960 375 13096 13065 24 25 12952 SDFFNSRXL $T=1361600 1517410 0 180 $X=1349640 $Y=1513470
X1347 12411 13061 13112 11960 375 13096 13186 24 25 13133 SDFFNSRXL $T=1351480 1517410 0 0 $X=1351478 $Y=1517158
X1348 12597 13149 13125 13102 337 12925 12827 24 25 13032 SDFFNSRXL $T=1363440 1473130 1 180 $X=1351480 $Y=1472878
X1349 12957 12795 13123 11960 337 12805 13146 24 25 13099 SDFFNSRXL $T=1352400 1554310 0 0 $X=1352398 $Y=1554058
X1350 366 13056 13126 13102 375 12926 13170 24 25 13109 SDFFNSRXL $T=1352860 1399330 1 0 $X=1352858 $Y=1395390
X1351 12597 12930 13138 13102 12641 12399 13149 24 25 13131 SDFFNSRXL $T=1354700 1465750 0 0 $X=1354698 $Y=1465498
X1352 13272 13258 13182 13102 375 13152 13027 24 25 13124 SDFFNSRXL $T=1367120 1443610 0 180 $X=1355160 $Y=1439670
X1353 289 13064 13154 379 380 12818 13240 24 25 395 SDFFNSRXL $T=1355620 1355050 0 0 $X=1355618 $Y=1354798
X1354 12942 13108 13155 13102 402 12688 13258 24 25 13260 SDFFNSRXL $T=1355620 1436230 1 0 $X=1355618 $Y=1432290
X1355 12597 370 13261 13102 381 12615 13055 24 25 13066 SDFFNSRXL $T=1367580 1480510 0 180 $X=1355620 $Y=1476570
X1356 12957 13139 13160 11960 402 13267 13279 24 25 13145 SDFFNSRXL $T=1356080 1569070 1 0 $X=1356078 $Y=1565130
X1357 366 13240 13136 379 380 12818 13117 24 25 13147 SDFFNSRXL $T=1368040 1362430 1 180 $X=1356080 $Y=1362178
X1358 13298 13270 13266 11960 13225 12692 13014 24 25 13129 SDFFNSRXL $T=1368040 1554310 0 180 $X=1356080 $Y=1550370
X1359 12957 13146 13134 11960 375 12805 13139 24 25 13118 SDFFNSRXL $T=1368040 1561690 1 180 $X=1356080 $Y=1561438
X1360 12942 13170 13174 13102 381 12462 13156 24 25 13158 SDFFNSRXL $T=1357920 1414090 1 0 $X=1357918 $Y=1410150
X1361 13298 13292 13287 11960 407 13042 13173 24 25 13165 SDFFNSRXL $T=1369880 1524790 1 180 $X=1357920 $Y=1524538
X1362 13294 13065 13303 13368 13225 12679 13419 24 25 13316 SDFFNSRXL $T=1368500 1502650 1 0 $X=1368498 $Y=1498710
X1363 366 13307 13311 13102 13225 12507 13367 24 25 13471 SDFFNSRXL $T=1369420 1391950 0 0 $X=1369418 $Y=1391698
X1364 13298 13173 13354 13368 431 13062 13376 24 25 13159 SDFFNSRXL $T=1370340 1532170 0 0 $X=1370338 $Y=1531918
X1365 366 13436 13319 13102 381 12683 13137 24 25 13318 SDFFNSRXL $T=1382760 1377190 1 180 $X=1370800 $Y=1376938
X1366 13294 13437 13423 13102 407 12560 13350 24 25 13315 SDFFNSRXL $T=1382760 1458370 1 180 $X=1370800 $Y=1458118
X1367 12957 13279 13435 13368 402 12805 13355 24 25 13317 SDFFNSRXL $T=1382760 1561690 1 180 $X=1370800 $Y=1561438
X1368 13272 13357 13364 13102 402 12508 13437 24 25 13424 SDFFNSRXL $T=1371260 1450990 0 0 $X=1371258 $Y=1450738
X1369 12942 13156 13361 13102 402 12462 13474 24 25 13488 SDFFNSRXL $T=1371720 1406710 0 0 $X=1371718 $Y=1406458
X1370 13294 13408 13442 13368 402 13025 13366 24 25 13353 SDFFNSRXL $T=1383680 1510030 1 180 $X=1371720 $Y=1509778
X1371 13272 13362 13381 13102 13225 12398 13385 24 25 13410 SDFFNSRXL $T=1372640 1428850 1 0 $X=1372638 $Y=1424910
X1372 13272 13385 13472 13102 407 13383 13369 24 25 13308 SDFFNSRXL $T=1384600 1428850 1 180 $X=1372640 $Y=1428598
X1373 13298 13409 13428 13368 13225 12692 13270 24 25 13310 SDFFNSRXL $T=1384600 1554310 0 180 $X=1372640 $Y=1550370
X1374 366 13380 13388 379 13225 12818 13440 24 25 13432 SDFFNSRXL $T=1373100 1362430 0 0 $X=1373098 $Y=1362178
X1375 12942 13481 13412 13102 13225 13391 13307 24 25 13282 SDFFNSRXL $T=1385060 1406710 0 180 $X=1373100 $Y=1402770
X1376 13272 13369 13478 13102 13225 12688 13382 24 25 13370 SDFFNSRXL $T=1385060 1436230 0 180 $X=1373100 $Y=1432290
X1377 12411 13483 13365 13368 402 12721 13292 24 25 13322 SDFFNSRXL $T=1385060 1524790 0 180 $X=1373100 $Y=1520850
X1378 13294 13419 13431 13368 402 13397 13387 24 25 13359 SDFFNSRXL $T=1385520 1495270 0 180 $X=1373560 $Y=1491330
X1379 12942 13474 13356 13102 13225 12687 13362 24 25 13244 SDFFNSRXL $T=1385980 1421470 0 180 $X=1374020 $Y=1417530
X1380 13294 13350 13438 13102 13225 12399 13395 24 25 13351 SDFFNSRXL $T=1385980 1465750 1 180 $X=1374020 $Y=1465498
X1381 12411 13366 13494 13368 13225 13096 13406 24 25 13305 SDFFNSRXL $T=1387360 1517410 1 180 $X=1375400 $Y=1517158
X1382 13294 13411 13439 13368 13225 13413 13408 24 25 13309 SDFFNSRXL $T=1387820 1502650 1 180 $X=1375860 $Y=1502398
X1383 13298 13376 13399 13368 431 12497 13409 24 25 13379 SDFFNSRXL $T=1387820 1539550 1 180 $X=1375860 $Y=1539298
X1384 13294 13387 13498 13368 431 12678 13411 24 25 13384 SDFFNSRXL $T=1388280 1487890 1 180 $X=1376320 $Y=1487638
X1385 366 430 13414 379 435 441 13380 24 25 445 SDFFNSRXL $T=1376780 1355050 0 0 $X=1376778 $Y=1354798
X1386 13294 13512 13504 13102 431 13425 13418 24 25 13396 SDFFNSRXL $T=1389660 1473130 1 180 $X=1377700 $Y=1472878
X1387 13294 13418 13441 13368 402 12615 13420 24 25 13373 SDFFNSRXL $T=1389660 1480510 1 180 $X=1377700 $Y=1480258
X1388 366 13509 13521 379 431 13475 437 24 25 13443 SDFFNSRXL $T=1393800 1369810 0 180 $X=1381840 $Y=1365870
X1389 13294 13513 13574 13368 447 12679 13479 24 25 13405 SDFFNSRXL $T=1394260 1495270 1 180 $X=1382300 $Y=1495018
X1390 12942 13580 13529 13102 381 13485 13477 24 25 13473 SDFFNSRXL $T=1394720 1391950 1 180 $X=1382760 $Y=1391698
X1391 13590 13510 13500 13368 447 12342 13483 24 25 13402 SDFFNSRXL $T=1395180 1532170 0 180 $X=1383220 $Y=1528230
X1392 13272 13491 13493 13102 447 12787 13357 24 25 13482 SDFFNSRXL $T=1384140 1443610 0 0 $X=1384138 $Y=1443358
X1393 13294 13492 13495 13102 402 12925 13512 24 25 13595 SDFFNSRXL $T=1384140 1473130 1 0 $X=1384138 $Y=1469190
X1394 13272 13496 13587 13102 431 13152 13491 24 25 13433 SDFFNSRXL $T=1396560 1443610 0 180 $X=1384600 $Y=1439670
X1395 13298 13355 13506 13368 402 13267 13575 24 25 13520 SDFFNSRXL $T=1385520 1561690 0 0 $X=1385518 $Y=1561438
X1396 13272 13382 13531 13102 402 13503 13496 24 25 13417 SDFFNSRXL $T=1397480 1421470 1 180 $X=1385520 $Y=1421218
X1397 13272 13585 13599 13102 431 12687 13501 24 25 13427 SDFFNSRXL $T=1397940 1421470 0 180 $X=1385980 $Y=1417530
X1398 13294 13420 13601 13368 431 13413 13499 24 25 13378 SDFFNSRXL $T=1397940 1502650 0 180 $X=1385980 $Y=1498710
X1399 13590 13406 13603 13368 407 13096 13502 24 25 13398 SDFFNSRXL $T=1397940 1517410 0 180 $X=1385980 $Y=1513470
X1400 12942 13484 13508 13102 407 13391 13525 24 25 13624 SDFFNSRXL $T=1386440 1406710 1 0 $X=1386438 $Y=1402770
X1401 13590 13606 13518 13368 447 13062 13510 24 25 13505 SDFFNSRXL $T=1398860 1532170 1 180 $X=1386900 $Y=1531918
X1402 366 13610 13579 379 431 12506 13509 24 25 13415 SDFFNSRXL $T=1399320 1377190 0 180 $X=1387360 $Y=1373250
X1403 13590 13536 13597 13368 447 12684 13513 24 25 13401 SDFFNSRXL $T=1399780 1510030 0 180 $X=1387820 $Y=1506090
X1404 13298 13514 13612 13368 431 12497 13519 24 25 13511 SDFFNSRXL $T=1399780 1539550 1 180 $X=1387820 $Y=1539298
X1405 13298 13616 13594 13368 13225 12692 13514 24 25 13507 SDFFNSRXL $T=1399780 1554310 0 180 $X=1387820 $Y=1550370
X1406 366 13440 13615 379 431 12818 13516 24 25 440 SDFFNSRXL $T=1400240 1362430 0 180 $X=1388280 $Y=1358490
X1407 13272 13593 13607 13102 453 12688 13523 24 25 13522 SDFFNSRXL $T=1401160 1436230 0 180 $X=1389200 $Y=1432290
X1408 13272 13501 13619 13102 447 13530 13526 24 25 13490 SDFFNSRXL $T=1401620 1414090 1 180 $X=1389660 $Y=1413838
X1409 12942 13525 13538 13102 13225 12462 13481 24 25 13613 SDFFNSRXL $T=1390580 1406710 0 0 $X=1390578 $Y=1406458
X1410 448 13534 13539 13368 454 13651 13654 24 25 13662 SDFFNSRXL $T=1390580 1480510 0 0 $X=1390578 $Y=1480258
X1411 13294 13533 13515 13102 407 12508 13532 24 25 13527 SDFFNSRXL $T=1402540 1450990 0 180 $X=1390580 $Y=1447050
X1412 13294 13654 13650 13102 454 13425 13492 24 25 13528 SDFFNSRXL $T=1402540 1480510 0 180 $X=1390580 $Y=1476570
X1413 13590 13582 13611 13368 431 13042 13536 24 25 13375 SDFFNSRXL $T=1402540 1524790 1 180 $X=1390580 $Y=1524538
X1414 366 13537 13573 13102 455 13655 13610 24 25 13665 SDFFNSRXL $T=1391040 1377190 0 0 $X=1391038 $Y=1376938
X1415 13298 13575 13578 13368 454 12805 13616 24 25 13670 SDFFNSRXL $T=1391500 1561690 1 0 $X=1391498 $Y=1557750
X1416 366 13516 13591 379 457 13475 13592 24 25 13617 SDFFNSRXL $T=1393800 1369810 1 0 $X=1393798 $Y=1365870
X1417 448 13479 13596 13368 455 12679 13678 24 25 13589 SDFFNSRXL $T=1394260 1495270 0 0 $X=1394258 $Y=1495018
X1418 13659 13677 13605 13102 431 12507 13580 24 25 13524 SDFFNSRXL $T=1406220 1391950 0 180 $X=1394260 $Y=1388010
X1419 366 13592 13598 379 455 441 456 24 25 460 SDFFNSRXL $T=1394720 1355050 1 0 $X=1394718 $Y=1351110
X1420 13590 13502 13583 13368 454 13096 13582 24 25 13623 SDFFNSRXL $T=1394720 1517410 0 0 $X=1394718 $Y=1517158
X1421 13294 13683 13622 13102 431 13576 13593 24 25 13588 SDFFNSRXL $T=1406680 1465750 0 180 $X=1394720 $Y=1461810
X1422 13272 13523 13581 13102 453 12398 13585 24 25 13716 SDFFNSRXL $T=1395180 1428850 1 0 $X=1395178 $Y=1424910
X1423 13272 13532 13653 13102 457 13152 13694 24 25 13656 SDFFNSRXL $T=1399780 1436230 0 0 $X=1399778 $Y=1435978
X1424 13590 13724 13675 13368 455 13062 13606 24 25 13652 SDFFNSRXL $T=1412660 1532170 1 180 $X=1400700 $Y=1531918
X1425 13659 13663 13666 13102 457 13476 13715 24 25 13758 SDFFNSRXL $T=1401620 1384570 0 0 $X=1401618 $Y=1384318
X1426 13298 13519 13667 13368 455 12497 13752 24 25 13756 SDFFNSRXL $T=1401620 1539550 0 0 $X=1401618 $Y=1539298
X1427 13704 13703 13719 13102 455 13668 13661 24 25 13614 SDFFNSRXL $T=1413580 1450990 1 180 $X=1401620 $Y=1450738
X1428 448 13672 13755 13368 13723 13651 13669 24 25 13577 SDFFNSRXL $T=1414960 1480510 1 180 $X=1403000 $Y=1480258
X1429 13294 13721 13684 13368 454 12678 13672 24 25 13657 SDFFNSRXL $T=1414960 1487890 1 180 $X=1403000 $Y=1487638
X1430 13659 13673 13681 13102 454 13485 13697 24 25 13771 SDFFNSRXL $T=1403460 1399330 1 0 $X=1403458 $Y=1395390
X1431 13590 13499 13682 13368 455 12684 13759 24 25 13761 SDFFNSRXL $T=1403460 1510030 1 0 $X=1403458 $Y=1506090
X1432 13789 13759 13757 13368 13723 13025 13676 24 25 13609 SDFFNSRXL $T=1415420 1510030 1 180 $X=1403460 $Y=1509778
X1433 470 13765 13760 379 13723 12506 13663 24 25 13604 SDFFNSRXL $T=1415880 1377190 0 180 $X=1403920 $Y=1373250
X1434 13590 13752 13692 13368 457 12974 13679 24 25 13618 SDFFNSRXL $T=1415880 1546930 0 180 $X=1403920 $Y=1542990
X1435 13590 13679 13763 13368 13723 12692 13680 24 25 13626 SDFFNSRXL $T=1415880 1554310 0 180 $X=1403920 $Y=1550370
X1436 13298 13680 13691 13368 454 12805 13764 24 25 13798 SDFFNSRXL $T=1404380 1561690 1 0 $X=1404378 $Y=1557750
X1437 13272 13690 13693 13102 454 13530 13707 24 25 13775 SDFFNSRXL $T=1404840 1414090 1 0 $X=1404838 $Y=1410150
X1438 366 13695 13700 379 457 13475 13765 24 25 13779 SDFFNSRXL $T=1405760 1369810 1 0 $X=1405758 $Y=1365870
X1439 13659 13773 13706 379 457 441 13695 24 25 459 SDFFNSRXL $T=1417720 1355050 1 180 $X=1405760 $Y=1354798
X1440 448 13678 13705 13368 454 13397 13721 24 25 13785 SDFFNSRXL $T=1406220 1495270 1 0 $X=1406218 $Y=1491330
X1441 13272 13526 13709 13102 455 13530 13777 24 25 13701 SDFFNSRXL $T=1406680 1414090 0 0 $X=1406678 $Y=1413838
X1442 13590 13699 13708 13368 454 13042 13724 24 25 13780 SDFFNSRXL $T=1406680 1524790 0 0 $X=1406678 $Y=1524538
X1443 13659 13697 13686 13102 457 13655 13537 24 25 13627 SDFFNSRXL $T=1418640 1377190 1 180 $X=1406680 $Y=1376938
X1444 13272 13707 13687 13102 13723 13391 13673 24 25 13753 SDFFNSRXL $T=1407140 1406710 1 0 $X=1407138 $Y=1402770
X1445 13704 13694 13751 13102 13723 12787 13703 24 25 13625 SDFFNSRXL $T=1419100 1443610 1 180 $X=1407140 $Y=1443358
X1446 13272 13784 13776 466 455 13485 13677 24 25 13702 SDFFNSRXL $T=1419560 1391950 1 180 $X=1407600 $Y=1391698
X1447 448 13696 13781 13766 13723 12925 13713 24 25 13608 SDFFNSRXL $T=1419560 1473130 0 180 $X=1407600 $Y=1469190
X1448 448 13713 13782 13766 457 13651 13534 24 25 13535 SDFFNSRXL $T=1419560 1487890 0 180 $X=1407600 $Y=1483950
X1449 13789 13676 13783 13368 457 12721 13711 24 25 13602 SDFFNSRXL $T=1419560 1517410 1 180 $X=1407600 $Y=1517158
X1450 13789 13711 13685 13368 454 12721 13699 24 25 13664 SDFFNSRXL $T=1419560 1524790 0 180 $X=1407600 $Y=1520850
X1451 13659 13715 13722 13102 13723 13476 13788 24 25 13787 SDFFNSRXL $T=1408060 1384570 1 0 $X=1408058 $Y=1380630
X1452 13704 13661 13720 13102 454 13576 13712 24 25 13791 SDFFNSRXL $T=1408060 1458370 0 0 $X=1408058 $Y=1458118
X1453 448 13669 13769 13766 457 13425 13683 24 25 13600 SDFFNSRXL $T=1420020 1473130 1 180 $X=1408060 $Y=1472878
X1454 13704 13777 13790 466 457 12687 13690 24 25 13671 SDFFNSRXL $T=1421400 1421470 0 180 $X=1409440 $Y=1417530
X1455 13704 13750 13710 13766 13723 12688 13714 24 25 13688 SDFFNSRXL $T=1421400 1436230 0 180 $X=1409440 $Y=1432290
X1456 13704 13832 13829 13766 454 13152 13750 24 25 13748 SDFFNSRXL $T=1423700 1436230 1 180 $X=1411740 $Y=1435978
X1457 13704 13689 13796 13766 13723 12398 13868 24 25 13895 SDFFNSRXL $T=1418640 1428850 1 0 $X=1418638 $Y=1424910
X1458 13789 13887 13884 13368 13723 13413 13792 24 25 13749 SDFFNSRXL $T=1430600 1502650 1 180 $X=1418640 $Y=1502398
X1459 448 13824 13828 13766 469 13425 13840 24 25 13896 SDFFNSRXL $T=1420480 1480510 1 0 $X=1420478 $Y=1476570
X1460 13272 13833 13898 466 13723 13391 13827 24 25 13767 SDFFNSRXL $T=1432900 1406710 0 180 $X=1420940 $Y=1402770
X1461 13928 13860 13897 13766 457 13576 13830 24 25 13754 SDFFNSRXL $T=1432900 1458370 1 180 $X=1420940 $Y=1458118
X1462 470 481 13825 466 473 441 13773 24 25 467 SDFFNSRXL $T=1433360 1355050 1 180 $X=1421400 $Y=1354798
X1463 448 13834 13841 13766 475 13651 13824 24 25 13925 SDFFNSRXL $T=1421860 1487890 1 0 $X=1421858 $Y=1483950
X1464 13659 13788 13838 466 447 13476 13862 24 25 13946 SDFFNSRXL $T=1422320 1384570 0 0 $X=1422318 $Y=1384318
X1465 13659 13839 13835 466 13723 13530 13833 24 25 13927 SDFFNSRXL $T=1422320 1414090 1 0 $X=1422318 $Y=1410150
X1466 448 13792 13883 13766 457 12679 13834 24 25 13725 SDFFNSRXL $T=1434280 1495270 1 180 $X=1422320 $Y=1495018
X1467 13789 13848 13843 13368 13723 12342 13837 24 25 13770 SDFFNSRXL $T=1434280 1532170 0 180 $X=1422320 $Y=1528230
X1468 13590 13764 13846 13368 454 12805 13842 24 25 13831 SDFFNSRXL $T=1422780 1554310 0 0 $X=1422778 $Y=1554058
X1469 13704 13830 13856 13766 13723 13668 13847 24 25 13768 SDFFNSRXL $T=1435200 1450990 1 180 $X=1423240 $Y=1450738
X1470 13659 13849 13859 466 477 13655 13882 24 25 13965 SDFFNSRXL $T=1423700 1377190 1 0 $X=1423698 $Y=1373250
X1471 13704 13851 13855 13766 478 13152 13832 24 25 13947 SDFFNSRXL $T=1423700 1436230 0 0 $X=1423698 $Y=1435978
X1472 13789 13857 13863 13368 469 13025 13881 24 25 13899 SDFFNSRXL $T=1424160 1510030 0 0 $X=1424158 $Y=1509778
X1473 13659 13862 13869 466 479 12507 13873 24 25 13952 SDFFNSRXL $T=1424620 1391950 1 0 $X=1424618 $Y=1388010
X1474 13659 13882 13931 466 478 13475 13858 24 25 13852 SDFFNSRXL $T=1436580 1369810 0 180 $X=1424620 $Y=1365870
X1475 13928 13935 13934 13766 480 13576 13860 24 25 13853 SDFFNSRXL $T=1436580 1465750 0 180 $X=1424620 $Y=1461810
X1476 13948 13870 13926 13368 475 12721 13857 24 25 13854 SDFFNSRXL $T=1436580 1517410 1 180 $X=1424620 $Y=1517158
X1477 13704 13868 13874 466 478 12687 13839 24 25 13976 SDFFNSRXL $T=1425080 1421470 1 0 $X=1425078 $Y=1417530
X1478 13948 13837 13938 13368 480 13042 13870 24 25 13861 SDFFNSRXL $T=1437040 1524790 1 180 $X=1425080 $Y=1524538
X1479 13948 13842 13936 13368 13723 12692 13866 24 25 13786 SDFFNSRXL $T=1437040 1554310 0 180 $X=1425080 $Y=1550370
X1480 13659 13873 13878 466 478 12926 13784 24 25 13953 SDFFNSRXL $T=1425540 1399330 0 0 $X=1425538 $Y=1399078
X1481 448 13840 13942 13766 482 13651 13875 24 25 13865 SDFFNSRXL $T=1437500 1480510 1 180 $X=1425540 $Y=1480258
X1482 13948 13866 13943 13368 457 12974 13872 24 25 13778 SDFFNSRXL $T=1437500 1546930 0 180 $X=1425540 $Y=1542990
X1483 13659 13858 13880 466 447 12818 13893 24 25 13989 SDFFNSRXL $T=1426000 1362430 0 0 $X=1425998 $Y=1362178
X1484 13948 13872 13944 13368 482 12497 13864 24 25 13871 SDFFNSRXL $T=1437960 1539550 0 180 $X=1426000 $Y=1535610
X1485 13789 14037 13967 13766 487 13413 13887 24 25 13929 SDFFNSRXL $T=1444400 1502650 1 180 $X=1432440 $Y=1502398
X1486 13948 13881 13956 13368 491 12721 13972 24 25 13970 SDFFNSRXL $T=1436580 1517410 0 0 $X=1436578 $Y=1517158
X1487 13659 13961 13968 466 480 12506 13849 24 25 14113 SDFFNSRXL $T=1437500 1369810 0 0 $X=1437498 $Y=1369558
X1488 13659 14068 13981 466 475 12683 13961 24 25 13950 SDFFNSRXL $T=1449460 1377190 1 180 $X=1437500 $Y=1376938
X1489 13704 13966 13963 13766 487 13383 13957 24 25 14149 SDFFNSRXL $T=1437960 1428850 0 0 $X=1437958 $Y=1428598
X1490 448 13875 13974 13766 487 13651 14042 24 25 13954 SDFFNSRXL $T=1437960 1487890 1 0 $X=1437958 $Y=1483950
X1491 13704 13973 13979 13766 480 12508 14061 24 25 13969 SDFFNSRXL $T=1438420 1450990 1 0 $X=1438418 $Y=1447050
X1492 13704 13957 14035 13766 482 13152 13973 24 25 13949 SDFFNSRXL $T=1450380 1436230 1 180 $X=1438420 $Y=1435978
X1493 13928 13992 14036 13766 493 12399 13935 24 25 13964 SDFFNSRXL $T=1450380 1465750 1 180 $X=1438420 $Y=1465498
X1494 13948 13990 13999 13368 480 12974 13997 24 25 14062 SDFFNSRXL $T=1439800 1546930 1 0 $X=1439798 $Y=1542990
X1495 13948 13997 14004 13368 469 12692 14047 24 25 14071 SDFFNSRXL $T=1440260 1554310 1 0 $X=1440258 $Y=1550370
X1496 13704 13984 14120 466 475 12687 13966 24 25 13983 SDFFNSRXL $T=1452220 1421470 0 180 $X=1440260 $Y=1417530
X1497 13789 14042 14003 13766 491 13397 13995 24 25 13993 SDFFNSRXL $T=1452680 1495270 0 180 $X=1440720 $Y=1491330
X1498 13659 14006 13975 466 469 13485 14002 24 25 14137 SDFFNSRXL $T=1441180 1399330 1 0 $X=1441178 $Y=1395390
X1499 13704 14130 13991 13766 480 13503 13984 24 25 13982 SDFFNSRXL $T=1453140 1421470 1 180 $X=1441180 $Y=1421218
X1500 13948 14046 14076 13368 475 12497 13990 24 25 14005 SDFFNSRXL $T=1453600 1539550 0 180 $X=1441640 $Y=1535610
X1501 13272 13827 14034 466 482 12462 14006 24 25 13962 SDFFNSRXL $T=1442100 1406710 0 0 $X=1442098 $Y=1406458
X1502 13948 13972 14048 13368 491 13042 14116 24 25 14115 SDFFNSRXL $T=1442100 1524790 0 0 $X=1442098 $Y=1524538
X1503 13789 14054 14132 13766 493 13397 14043 24 25 13985 SDFFNSRXL $T=1454060 1487890 1 180 $X=1442100 $Y=1487638
X1504 13789 14116 14055 13766 496 12684 14037 24 25 14031 SDFFNSRXL $T=1454060 1510030 0 180 $X=1442100 $Y=1506090
X1505 13948 14140 14136 13368 487 12342 14046 24 25 14038 SDFFNSRXL $T=1454520 1532170 0 180 $X=1442560 $Y=1528230
X1506 13928 14049 13977 13766 491 12560 13992 24 25 14152 SDFFNSRXL $T=1443020 1458370 1 0 $X=1443018 $Y=1454430
X1507 13789 14043 14143 13766 496 13425 14051 24 25 13940 SDFFNSRXL $T=1455440 1480510 0 180 $X=1443480 $Y=1476570
X1508 13789 13995 14121 13766 496 12679 14054 24 25 13971 SDFFNSRXL $T=1456360 1495270 1 180 $X=1444400 $Y=1495018
X1509 13704 14061 14069 13766 487 13668 14049 24 25 14184 SDFFNSRXL $T=1446700 1450990 0 0 $X=1446698 $Y=1450738
X1510 14194 14181 14229 13766 502 13025 14123 24 25 14070 SDFFNSRXL $T=1462340 1510030 1 180 $X=1450380 $Y=1509778
X1511 13659 14128 14129 466 494 12506 14041 24 25 14239 SDFFNSRXL $T=1450840 1369810 0 0 $X=1450838 $Y=1369558
X1512 13928 14148 14156 466 493 12507 14157 24 25 14179 SDFFNSRXL $T=1453600 1391950 1 0 $X=1453598 $Y=1388010
X1513 13659 14157 14167 466 504 12683 14068 24 25 14244 SDFFNSRXL $T=1454980 1377190 0 0 $X=1454978 $Y=1376938
X1514 13789 14051 14169 13766 14228 12678 14268 24 25 14227 SDFFNSRXL $T=1454980 1487890 1 0 $X=1454978 $Y=1483950
X1515 14158 14166 14172 13766 496 13576 14265 24 25 14248 SDFFNSRXL $T=1455440 1465750 1 0 $X=1455438 $Y=1461810
X1516 14158 14235 14064 13766 491 13152 14119 24 25 14159 SDFFNSRXL $T=1467400 1443610 0 180 $X=1455440 $Y=1439670
X1517 14158 14265 14238 13766 504 12399 14164 24 25 14160 SDFFNSRXL $T=1467400 1465750 1 180 $X=1455440 $Y=1465498
X1518 14158 14164 14174 13766 14228 12560 14267 24 25 14272 SDFFNSRXL $T=1455900 1458370 1 0 $X=1455898 $Y=1454430
X1519 14282 14233 14171 13766 493 13383 14130 24 25 14163 SDFFNSRXL $T=1467860 1428850 1 180 $X=1455900 $Y=1428598
X1520 13789 14268 14245 13766 504 13397 14176 24 25 14175 SDFFNSRXL $T=1469240 1487890 1 180 $X=1457280 $Y=1487638
X1521 14194 14243 14277 14256 14228 12342 14140 24 25 14178 SDFFNSRXL $T=1469700 1532170 0 180 $X=1457740 $Y=1528230
X1522 14194 14190 14278 14256 482 12974 14186 24 25 14180 SDFFNSRXL $T=1470160 1546930 0 180 $X=1458200 $Y=1542990
X1523 470 13994 14225 466 504 441 513 24 25 14266 SDFFNSRXL $T=1458660 1355050 0 0 $X=1458658 $Y=1354798
X1524 14158 14119 14234 13766 496 13152 14317 24 25 14262 SDFFNSRXL $T=1459120 1436230 0 0 $X=1459118 $Y=1435978
X1525 14194 14047 14191 14256 469 12805 14190 24 25 14250 SDFFNSRXL $T=1459120 1554310 1 0 $X=1459118 $Y=1550370
X1526 13928 14188 14231 466 482 12926 14148 24 25 14195 SDFFNSRXL $T=1459580 1399330 1 0 $X=1459578 $Y=1395390
X1527 14194 14176 14189 13766 504 13413 14181 24 25 14193 SDFFNSRXL $T=1459580 1502650 1 0 $X=1459578 $Y=1498710
X1528 14158 14267 14283 13766 493 13668 14235 24 25 14192 SDFFNSRXL $T=1471540 1450990 1 180 $X=1459580 $Y=1450738
X1529 14194 14186 14284 14256 482 12974 14236 24 25 14053 SDFFNSRXL $T=1471540 1546930 1 180 $X=1459580 $Y=1546678
X1530 13928 14138 14170 466 496 12926 14188 24 25 14279 SDFFNSRXL $T=1460040 1399330 0 0 $X=1460038 $Y=1399078
X1531 14282 14321 14275 13766 504 13503 14233 24 25 14226 SDFFNSRXL $T=1472000 1421470 1 180 $X=1460040 $Y=1421218
X1532 14194 14123 14260 13766 14228 13025 14274 24 25 14254 SDFFNSRXL $T=1462340 1510030 0 0 $X=1462338 $Y=1509778
X1533 14158 14259 14330 13766 14228 12925 14249 24 25 14242 SDFFNSRXL $T=1474300 1473130 0 180 $X=1462340 $Y=1469190
X1534 470 508 14261 466 493 12506 14340 24 25 14338 SDFFNSRXL $T=1462800 1369810 0 0 $X=1462798 $Y=1369558
X1535 14158 14331 14333 13766 14228 13425 14259 24 25 14246 SDFFNSRXL $T=1474760 1473130 1 180 $X=1462800 $Y=1472878
X1536 14194 14274 14341 14256 14228 13096 14263 24 25 14251 SDFFNSRXL $T=1475680 1517410 0 180 $X=1463720 $Y=1513470
X1537 14282 14313 14320 466 480 12462 14379 24 25 14413 SDFFNSRXL $T=1469240 1406710 0 0 $X=1469238 $Y=1406458
X1538 13789 14315 14322 13766 496 13397 14331 24 25 14378 SDFFNSRXL $T=1469240 1487890 0 0 $X=1469238 $Y=1487638
X1539 14282 14319 14323 466 469 13391 14313 24 25 14416 SDFFNSRXL $T=1469700 1406710 1 0 $X=1469698 $Y=1402770
X1540 14282 14379 14346 14370 504 13503 14328 24 25 14232 SDFFNSRXL $T=1483500 1421470 0 180 $X=1471540 $Y=1417530
X1541 14158 14375 14419 14370 14228 13668 14329 24 25 14325 SDFFNSRXL $T=1483960 1450990 1 180 $X=1472000 $Y=1450738
X1542 14194 14352 14360 14256 480 12497 14332 24 25 14237 SDFFNSRXL $T=1483960 1539550 0 180 $X=1472000 $Y=1535610
X1543 470 518 14422 466 482 12818 14334 24 25 14326 SDFFNSRXL $T=1484420 1355050 1 180 $X=1472460 $Y=1354798
X1544 14282 14345 14350 466 504 13476 14128 24 25 14271 SDFFNSRXL $T=1484420 1384570 1 180 $X=1472460 $Y=1384318
X1545 14282 14359 14336 14370 14228 13503 14321 24 25 14314 SDFFNSRXL $T=1484420 1421470 1 180 $X=1472460 $Y=1421218
X1546 13789 14339 14343 13766 487 12679 14315 24 25 14411 SDFFNSRXL $T=1472920 1495270 1 0 $X=1472918 $Y=1491330
X1547 14282 14427 14425 466 479 13391 14319 24 25 14335 SDFFNSRXL $T=1484880 1399330 1 180 $X=1472920 $Y=1399078
X1548 14158 14412 14426 14370 480 12399 14166 24 25 14337 SDFFNSRXL $T=1484880 1465750 0 180 $X=1472920 $Y=1461810
X1549 14158 14317 14347 13766 469 13152 14375 24 25 14517 SDFFNSRXL $T=1473380 1443610 1 0 $X=1473378 $Y=1439670
X1550 14282 14355 14429 466 504 13485 14345 24 25 14316 SDFFNSRXL $T=1485340 1391950 1 180 $X=1473380 $Y=1391698
X1551 14194 14380 14344 13766 519 13413 14339 24 25 14196 SDFFNSRXL $T=1485340 1502650 1 180 $X=1473380 $Y=1502398
X1552 14194 14263 14342 14256 519 13042 14252 24 25 14177 SDFFNSRXL $T=1485340 1524790 0 180 $X=1473380 $Y=1520850
X1553 14446 14249 14434 13766 519 12925 14348 24 25 14173 SDFFNSRXL $T=1486260 1473130 0 180 $X=1474300 $Y=1469190
X1554 470 14377 14435 466 496 12506 14349 24 25 14257 SDFFNSRXL $T=1486720 1369810 1 180 $X=1474760 $Y=1369558
X1555 14194 14443 14439 14256 475 12974 14352 24 25 14264 SDFFNSRXL $T=1487180 1546930 0 180 $X=1475220 $Y=1542990
X1556 14282 14340 14428 466 521 12683 14355 24 25 14327 SDFFNSRXL $T=1488100 1377190 1 180 $X=1476140 $Y=1376938
X1557 14158 14361 14367 14370 480 12688 14451 24 25 14458 SDFFNSRXL $T=1476600 1436230 1 0 $X=1476598 $Y=1432290
X1558 14158 14362 14364 14370 469 13576 14412 24 25 14465 SDFFNSRXL $T=1476600 1458370 0 0 $X=1476598 $Y=1458118
X1559 13789 14348 14365 13766 502 13651 14438 24 25 14423 SDFFNSRXL $T=1476600 1480510 0 0 $X=1476598 $Y=1480258
X1560 14194 14332 14368 14256 480 13062 14455 24 25 14440 SDFFNSRXL $T=1476600 1532170 1 0 $X=1476598 $Y=1528230
X1561 14282 14451 14444 14370 14228 12398 14359 24 25 14258 SDFFNSRXL $T=1488560 1428850 0 180 $X=1476600 $Y=1424910
X1562 14194 14236 14373 14256 469 12692 14443 24 25 14460 SDFFNSRXL $T=1477060 1546930 0 0 $X=1477058 $Y=1546678
X1563 14158 14371 14430 14370 504 12787 14361 24 25 14276 SDFFNSRXL $T=1489020 1443610 1 180 $X=1477060 $Y=1443358
X1564 14282 14328 14374 466 479 13530 14449 24 25 14414 SDFFNSRXL $T=1477520 1414090 0 0 $X=1477518 $Y=1413838
X1565 14194 14351 14372 14256 519 13025 14380 24 25 14471 SDFFNSRXL $T=1477520 1510030 0 0 $X=1477518 $Y=1509778
X1566 14158 14329 14436 14370 504 12508 14371 24 25 14269 SDFFNSRXL $T=1489480 1450990 0 180 $X=1477520 $Y=1447050
X1567 470 14334 14437 466 524 12818 14377 24 25 14281 SDFFNSRXL $T=1490400 1362430 1 180 $X=1478440 $Y=1362178
X1568 14194 14431 14353 14256 14228 12684 14351 24 25 14534 SDFFNSRXL $T=1483040 1510030 1 0 $X=1483038 $Y=1506090
X1569 14446 14438 14519 13766 491 12678 14447 24 25 14432 SDFFNSRXL $T=1497300 1487890 0 180 $X=1485340 $Y=1483950
X1570 14158 14525 14518 14370 475 12560 14362 24 25 14445 SDFFNSRXL $T=1497760 1458370 0 180 $X=1485800 $Y=1454430
X1571 14282 14513 14556 14370 479 13383 14457 24 25 14452 SDFFNSRXL $T=1499140 1428850 1 180 $X=1487180 $Y=1428598
X1572 14446 14447 14463 13766 487 12925 14536 24 25 14583 SDFFNSRXL $T=1488100 1473130 1 0 $X=1488098 $Y=1469190
X1573 14282 14468 14472 14370 487 13530 14513 24 25 14558 SDFFNSRXL $T=1489480 1414090 1 0 $X=1489478 $Y=1410150
X1574 14282 14449 14470 14370 475 12687 14468 24 25 14448 SDFFNSRXL $T=1489480 1414090 0 0 $X=1489478 $Y=1413838
X1575 14194 14455 14473 14256 487 13062 14526 24 25 14541 SDFFNSRXL $T=1489480 1532170 1 0 $X=1489478 $Y=1528230
X1576 14282 14551 14531 14370 480 12926 14427 24 25 14456 SDFFNSRXL $T=1501440 1399330 0 180 $X=1489480 $Y=1395390
X1577 470 14349 14511 530 504 13655 14537 24 25 14575 SDFFNSRXL $T=1489940 1369810 0 0 $X=1489938 $Y=1369558
X1578 14158 14515 14619 14370 479 12508 14525 24 25 14461 SDFFNSRXL $T=1504660 1450990 0 180 $X=1492700 $Y=1447050
X1579 14446 14536 14544 14256 496 13425 14640 24 25 14655 SDFFNSRXL $T=1493620 1480510 1 0 $X=1493618 $Y=1476570
X1580 470 14537 14548 530 487 12683 14567 24 25 14658 SDFFNSRXL $T=1494080 1377190 0 0 $X=1494078 $Y=1376938
X1581 14194 14542 14549 14256 480 12974 14532 24 25 14590 SDFFNSRXL $T=1494080 1539550 0 0 $X=1494078 $Y=1539298
X1582 14282 14638 14629 14370 475 13485 14543 24 25 14512 SDFFNSRXL $T=1506040 1391950 1 180 $X=1494080 $Y=1391698
X1583 14446 14526 14634 14256 482 13042 14542 24 25 14453 SDFFNSRXL $T=1506040 1524790 1 180 $X=1494080 $Y=1524538
X1584 14282 14457 14555 14370 496 13503 14554 24 25 14568 SDFFNSRXL $T=1494540 1421470 0 0 $X=1494538 $Y=1421218
X1585 14194 14532 14550 14256 482 12692 14647 24 25 14642 SDFFNSRXL $T=1494540 1546930 0 0 $X=1494538 $Y=1546678
X1586 14282 14543 14639 14370 495 13391 14551 24 25 14539 SDFFNSRXL $T=1506500 1399330 1 180 $X=1494540 $Y=1399078
X1587 14446 14564 14620 14256 496 13096 14431 24 25 14522 SDFFNSRXL $T=1506500 1510030 1 180 $X=1494540 $Y=1509778
X1588 14158 14585 14514 14370 475 12787 14515 24 25 14529 SDFFNSRXL $T=1506960 1443610 0 180 $X=1495000 $Y=1439670
X1589 14446 14570 14654 14256 504 13413 14564 24 25 14520 SDFFNSRXL $T=1508340 1502650 0 180 $X=1496380 $Y=1498710
X1590 531 14567 14573 530 495 13655 14668 24 25 14644 SDFFNSRXL $T=1496840 1377190 1 0 $X=1496838 $Y=1373250
X1591 14446 14667 14660 14256 487 12678 14570 24 25 14563 SDFFNSRXL $T=1509260 1487890 0 180 $X=1497300 $Y=1483950
X1592 531 14688 14553 530 496 12818 534 24 25 14581 SDFFNSRXL $T=1511560 1355050 1 180 $X=1499600 $Y=1354798
X1593 14158 14698 14586 14370 487 12787 14585 24 25 14579 SDFFNSRXL $T=1512480 1443610 1 180 $X=1500520 $Y=1443358
X1594 14657 14640 14675 14256 491 13425 14732 24 25 14617 SDFFNSRXL $T=1506960 1473130 0 0 $X=1506958 $Y=1472878
X1595 14770 14731 14662 14370 502 13485 14638 24 25 14656 SDFFNSRXL $T=1518920 1391950 1 180 $X=1506960 $Y=1391698
X1596 14446 14665 14691 14256 496 13025 14664 24 25 14653 SDFFNSRXL $T=1518920 1502650 1 180 $X=1506960 $Y=1502398
X1597 14446 14684 14758 14256 502 13025 14665 24 25 14560 SDFFNSRXL $T=1518920 1510030 0 180 $X=1506960 $Y=1506090
X1598 14158 14732 14677 14370 502 13668 14670 24 25 14621 SDFFNSRXL $T=1519380 1450990 1 180 $X=1507420 $Y=1450738
X1599 14659 14674 14682 14370 539 12787 14698 24 25 14768 SDFFNSRXL $T=1507880 1443610 1 0 $X=1507878 $Y=1439670
X1600 14659 14746 14761 14370 14228 13383 14674 24 25 14669 SDFFNSRXL $T=1519840 1428850 1 180 $X=1507880 $Y=1428598
X1601 14657 14767 14762 14370 502 12925 14678 24 25 14628 SDFFNSRXL $T=1519840 1465750 0 180 $X=1507880 $Y=1461810
X1602 14659 14649 14690 14370 14228 13503 14692 24 25 14776 SDFFNSRXL $T=1508800 1421470 1 0 $X=1508798 $Y=1417530
X1603 531 14668 14695 530 524 13655 14736 24 25 14775 SDFFNSRXL $T=1509260 1377190 1 0 $X=1509258 $Y=1373250
X1604 14659 14692 14766 14370 491 13530 14689 24 25 14523 SDFFNSRXL $T=1521220 1414090 0 180 $X=1509260 $Y=1410150
X1605 14657 14687 14772 14256 519 13425 14686 24 25 14671 SDFFNSRXL $T=1521220 1480510 0 180 $X=1509260 $Y=1476570
X1606 14657 14739 14773 14256 502 12678 14687 24 25 14546 SDFFNSRXL $T=1521220 1487890 0 180 $X=1509260 $Y=1483950
X1607 14657 14774 14740 14256 491 12679 14667 24 25 14530 SDFFNSRXL $T=1521220 1495270 0 180 $X=1509260 $Y=1491330
X1608 14446 14664 14699 14256 14228 13413 14774 24 25 14777 SDFFNSRXL $T=1509720 1495270 0 0 $X=1509718 $Y=1495018
X1609 13948 14733 14771 14256 491 13062 14729 24 25 14571 SDFFNSRXL $T=1522140 1524790 1 180 $X=1510180 $Y=1524538
X1610 13948 14647 14700 14256 475 12974 14741 24 25 14566 SDFFNSRXL $T=1510640 1539550 0 0 $X=1510638 $Y=1539298
X1611 14770 14751 14685 14370 491 12926 14731 24 25 14697 SDFFNSRXL $T=1523060 1399330 0 180 $X=1511100 $Y=1395390
X1612 14659 14670 14789 14370 491 13668 14735 24 25 14631 SDFFNSRXL $T=1523060 1450990 0 180 $X=1511100 $Y=1447050
X1613 531 14736 14742 530 453 13655 14821 24 25 14839 SDFFNSRXL $T=1511560 1369810 1 0 $X=1511558 $Y=1365870
X1614 531 538 14730 530 524 13475 14688 24 25 14635 SDFFNSRXL $T=1523520 1362430 1 180 $X=1511560 $Y=1362178
X1615 13948 14741 14694 14256 475 13062 14733 24 25 14420 SDFFNSRXL $T=1512020 1532170 0 0 $X=1512018 $Y=1531918
X1616 14657 14678 14784 14256 14228 12925 14739 24 25 14728 SDFFNSRXL $T=1523980 1473130 0 180 $X=1512020 $Y=1469190
X1617 14657 14747 14750 14370 14228 13576 14767 24 25 14743 SDFFNSRXL $T=1513400 1458370 0 0 $X=1513398 $Y=1458118
X1618 531 14840 14783 530 539 13476 14751 24 25 14748 SDFFNSRXL $T=1526280 1384570 1 180 $X=1514320 $Y=1384318
X1619 14446 14843 14785 14256 14228 13096 14693 24 25 14557 SDFFNSRXL $T=1526740 1510030 1 180 $X=1514780 $Y=1509778
X1620 14657 14735 14845 14370 539 13576 14747 24 25 14683 SDFFNSRXL $T=1527200 1458370 0 180 $X=1515240 $Y=1454430
X1621 14659 14760 14738 14370 519 13383 14746 24 25 14757 SDFFNSRXL $T=1517080 1428850 1 0 $X=1517078 $Y=1424910
X1622 14657 14930 14878 14256 544 12925 14836 24 25 14833 SDFFNSRXL $T=1535940 1473130 0 180 $X=1523980 $Y=1469190
X1623 13948 14676 14926 14256 519 13042 14837 24 25 14759 SDFFNSRXL $T=1535940 1524790 0 180 $X=1523980 $Y=1520850
X1624 14659 14929 14928 14370 519 13530 14842 24 25 14754 SDFFNSRXL $T=1536400 1414090 0 180 $X=1524440 $Y=1410150
X1625 13948 14729 14673 14256 14228 13062 14676 24 25 14782 SDFFNSRXL $T=1536400 1532170 0 180 $X=1524440 $Y=1528230
X1626 14770 14863 14933 14370 539 13391 14848 24 25 14763 SDFFNSRXL $T=1536860 1399330 1 180 $X=1524900 $Y=1399078
X1627 531 14852 14855 530 524 13475 14880 24 25 550 SDFFNSRXL $T=1526280 1355050 0 0 $X=1526278 $Y=1354798
X1628 14659 14952 14939 14370 544 13383 14853 24 25 14849 SDFFNSRXL $T=1538240 1421470 1 180 $X=1526280 $Y=1421218
X1629 14770 14848 14867 530 524 13485 14871 24 25 14820 SDFFNSRXL $T=1527200 1391950 1 0 $X=1527198 $Y=1388010
X1630 14657 14686 14868 14256 544 13651 14930 24 25 14971 SDFFNSRXL $T=1527200 1480510 1 0 $X=1527198 $Y=1476570
X1631 14657 14858 14841 14256 544 13397 14834 24 25 14982 SDFFNSRXL $T=1527200 1487890 1 0 $X=1527198 $Y=1483950
X1632 14446 14860 14953 14256 539 13025 14843 24 25 14769 SDFFNSRXL $T=1539160 1510030 0 180 $X=1527200 $Y=1506090
X1633 14659 14842 14864 14370 524 13391 14863 24 25 14823 SDFFNSRXL $T=1539620 1406710 0 180 $X=1527660 $Y=1402770
X1634 14446 14834 14875 14256 519 13397 14976 24 25 14755 SDFFNSRXL $T=1528580 1487890 0 0 $X=1528578 $Y=1487638
X1635 14446 14873 14850 14256 539 13413 14860 24 25 14764 SDFFNSRXL $T=1528580 1502650 1 0 $X=1528578 $Y=1498710
X1636 14770 14871 14927 530 519 13476 14840 24 25 14753 SDFFNSRXL $T=1541460 1384570 1 180 $X=1529500 $Y=1384318
X1637 568 15090 15081 14370 544 13668 14973 24 25 14915 SDFFNSRXL $T=1550660 1443610 1 180 $X=1538700 $Y=1443358
X1638 14657 14986 15034 14256 544 13397 15059 24 25 14981 SDFFNSRXL $T=1541460 1487890 0 0 $X=1541458 $Y=1487638
X1639 568 15138 15065 14370 519 13503 14952 24 25 14989 SDFFNSRXL $T=1553880 1421470 0 180 $X=1541920 $Y=1417530
X1640 14657 14973 15135 14370 544 13152 15031 24 25 14917 SDFFNSRXL $T=1553880 1436230 0 180 $X=1541920 $Y=1432290
X1641 565 15046 15055 530 453 13475 558 24 25 15030 SDFFNSRXL $T=1554340 1362430 0 180 $X=1542380 $Y=1358490
X1642 14657 14976 15053 14256 544 13413 15153 24 25 15035 SDFFNSRXL $T=1543760 1495270 1 0 $X=1543758 $Y=1491330
X1643 565 15155 15151 530 453 13655 15056 24 25 15046 SDFFNSRXL $T=1556640 1369810 0 180 $X=1544680 $Y=1365870
X1644 565 566 567 530 516 441 14922 24 25 571 SDFFNSRXL $T=1545600 1355050 1 0 $X=1545598 $Y=1351110
X1645 14659 15068 15071 14370 544 13391 15149 24 25 15051 SDFFNSRXL $T=1545600 1399330 1 0 $X=1545598 $Y=1395390
X1646 14659 15031 15072 14370 544 13383 15139 24 25 15039 SDFFNSRXL $T=1545600 1428850 1 0 $X=1545598 $Y=1424910
X1647 565 14880 15077 530 516 13475 14935 24 25 15188 SDFFNSRXL $T=1546060 1355050 0 0 $X=1546058 $Y=1354798
X1648 14657 15057 15078 14256 544 13651 15045 24 25 15166 SDFFNSRXL $T=1546060 1480510 0 0 $X=1546058 $Y=1480258
X1649 14657 15059 15058 14256 544 13397 15057 24 25 14969 SDFFNSRXL $T=1558020 1487890 0 180 $X=1546060 $Y=1483950
X1650 14659 15149 15044 14370 519 13485 15064 24 25 15066 SDFFNSRXL $T=1558480 1391950 1 180 $X=1546520 $Y=1391698
X1651 14657 15132 15136 14370 544 13668 15228 24 25 15164 SDFFNSRXL $T=1550660 1443610 0 0 $X=1550658 $Y=1443358
X1652 568 15267 15271 14370 544 13530 15176 24 25 15174 SDFFNSRXL $T=1570440 1414090 0 180 $X=1558480 $Y=1410150
X1653 14657 15231 15237 14256 544 13425 15253 24 25 15266 SDFFNSRXL $T=1560780 1473130 1 0 $X=1560778 $Y=1469190
X1654 565 15283 15246 586 453 13655 14925 24 25 15155 SDFFNSRXL $T=1573660 1369810 1 180 $X=1561700 $Y=1369558
X1655 565 15286 15282 586 453 13475 15242 24 25 15234 SDFFNSRXL $T=1574120 1362430 0 180 $X=1562160 $Y=1358490
X1656 14657 15240 15250 14256 544 13651 15231 24 25 15327 SDFFNSRXL $T=1563080 1480510 0 0 $X=1563078 $Y=1480258
X1657 565 15243 15254 586 453 13655 15187 24 25 15283 SDFFNSRXL $T=1563540 1377190 1 0 $X=1563538 $Y=1373250
X1658 568 15320 15328 14370 544 13530 15248 24 25 15185 SDFFNSRXL $T=1575500 1406710 0 180 $X=1563540 $Y=1402770
X1659 14659 585 15258 14370 519 13485 15334 24 25 15335 SDFFNSRXL $T=1564000 1391950 0 0 $X=1563998 $Y=1391698
X1660 568 15248 15256 14370 519 13503 15267 24 25 15284 SDFFNSRXL $T=1564000 1414090 0 0 $X=1563998 $Y=1413838
X1661 568 15249 15259 14370 544 13668 15324 24 25 15132 SDFFNSRXL $T=1564000 1450990 0 0 $X=1563998 $Y=1450738
X1662 14657 15253 15257 14370 544 13576 15249 24 25 15280 SDFFNSRXL $T=1564000 1458370 0 0 $X=1563998 $Y=1458118
X1663 565 15318 15239 586 544 13476 15243 24 25 15189 SDFFNSRXL $T=1576420 1377190 1 180 $X=1564460 $Y=1376938
X1664 14659 15244 15264 586 519 13476 15318 24 25 15323 SDFFNSRXL $T=1565380 1384570 0 0 $X=1565378 $Y=1384318
X1665 565 15188 15349 586 516 13475 15270 24 25 15286 SDFFNSRXL $T=1582860 1355050 1 180 $X=1570900 $Y=1354798
X1666 10157 25 10182 96 24 NOR2X1 $T=1129300 1362430 0 0 $X=1129298 $Y=1362178
X1667 10396 25 9920 10471 24 NOR2X1 $T=1148160 1450990 0 180 $X=1146780 $Y=1447050
X1668 10178 25 10065 10499 24 NOR2X1 $T=1155520 1355050 1 0 $X=1155518 $Y=1351110
X1669 10492 25 10467 10463 24 NOR2X1 $T=1157360 1480510 1 0 $X=1157358 $Y=1476570
X1670 10615 25 10599 10387 24 NOR2X1 $T=1163340 1517410 0 180 $X=1161960 $Y=1513470
X1671 118 25 131 10668 24 NOR2X1 $T=1164260 1355050 1 0 $X=1164258 $Y=1351110
X1672 10652 25 10628 10743 24 NOR2X1 $T=1170700 1458370 1 0 $X=1170698 $Y=1454430
X1673 10658 25 10628 10751 24 NOR2X1 $T=1171160 1391950 0 0 $X=1171158 $Y=1391698
X1674 10619 25 10628 10778 24 NOR2X1 $T=1172540 1391950 1 0 $X=1172538 $Y=1388010
X1675 10675 25 131 10806 24 NOR2X1 $T=1173000 1369810 1 0 $X=1172998 $Y=1365870
X1676 10607 25 10628 10797 24 NOR2X1 $T=1173920 1369810 0 0 $X=1173918 $Y=1369558
X1677 10656 25 10628 10767 24 NOR2X1 $T=1173920 1384570 0 0 $X=1173918 $Y=1384318
X1678 10618 25 10628 10800 24 NOR2X1 $T=1174380 1384570 1 0 $X=1174378 $Y=1380630
X1679 10712 25 10628 10768 24 NOR2X1 $T=1174380 1465750 1 0 $X=1174378 $Y=1461810
X1680 148 25 10806 10814 24 NOR2X1 $T=1178520 1377190 1 0 $X=1178518 $Y=1373250
X1681 10714 25 10628 10849 24 NOR2X1 $T=1178520 1436230 0 0 $X=1178518 $Y=1435978
X1682 10753 25 10628 10850 24 NOR2X1 $T=1178980 1473130 0 0 $X=1178978 $Y=1472878
X1683 150 25 10800 10861 24 NOR2X1 $T=1180360 1384570 0 180 $X=1178980 $Y=1380630
X1684 10774 25 10628 10863 24 NOR2X1 $T=1179900 1465750 0 0 $X=1179898 $Y=1465498
X1685 10925 25 155 11015 24 NOR2X1 $T=1185880 1355050 0 0 $X=1185878 $Y=1354798
X1686 10814 25 10861 11014 24 NOR2X1 $T=1187260 1377190 1 0 $X=1187258 $Y=1373250
X1687 10856 25 10628 11051 24 NOR2X1 $T=1190020 1443610 1 0 $X=1190018 $Y=1439670
X1688 11019 25 10628 11063 24 NOR2X1 $T=1191860 1465750 0 0 $X=1191858 $Y=1465498
X1689 10483 25 10628 11093 24 NOR2X1 $T=1193240 1465750 1 0 $X=1193238 $Y=1461810
X1690 11077 25 11015 171 24 NOR2X1 $T=1197840 1355050 0 180 $X=1196460 $Y=1351110
X1691 11123 25 10396 10615 24 NOR2X1 $T=1197840 1502650 0 180 $X=1196460 $Y=1498710
X1692 10908 25 11086 11172 24 NOR2X1 $T=1197380 1384570 1 0 $X=1197378 $Y=1380630
X1693 178 25 10668 11077 24 NOR2X1 $T=1205200 1355050 1 0 $X=1205198 $Y=1351110
X1694 176 25 10797 11297 24 NOR2X1 $T=1208880 1369810 1 0 $X=1208878 $Y=1365870
X1695 191 25 10767 11331 24 NOR2X1 $T=1213940 1377190 0 0 $X=1213938 $Y=1376938
X1696 11297 25 11331 11236 24 NOR2X1 $T=1214400 1377190 1 0 $X=1214398 $Y=1373250
X1697 11325 25 11332 11312 24 NOR2X1 $T=1214400 1384570 0 0 $X=1214398 $Y=1384318
X1698 11304 25 11472 11454 24 NOR2X1 $T=1224060 1399330 1 0 $X=1224058 $Y=1395390
X1699 11486 25 10778 11520 24 NOR2X1 $T=1225900 1384570 0 0 $X=1225898 $Y=1384318
X1700 11364 25 11051 11497 24 NOR2X1 $T=1227740 1443610 1 180 $X=1226360 $Y=1443358
X1701 11497 25 11502 11482 24 NOR2X1 $T=1226820 1436230 0 0 $X=1226818 $Y=1435978
X1702 11496 25 10751 11527 24 NOR2X1 $T=1227280 1399330 1 0 $X=1227278 $Y=1395390
X1703 11463 25 11063 11535 24 NOR2X1 $T=1231880 1480510 0 180 $X=1230500 $Y=1476570
X1704 11520 25 11527 11513 24 NOR2X1 $T=1230960 1391950 0 0 $X=1230958 $Y=1391698
X1705 11472 25 11543 11526 24 NOR2X1 $T=1230960 1406710 1 0 $X=1230958 $Y=1402770
X1706 11530 25 10849 11502 24 NOR2X1 $T=1231880 1436230 0 0 $X=1231878 $Y=1435978
X1707 11662 25 10736 11678 24 NOR2X1 $T=1239240 1369810 1 0 $X=1239238 $Y=1365870
X1708 11535 25 11673 11689 24 NOR2X1 $T=1239240 1473130 1 0 $X=1239238 $Y=1469190
X1709 11620 25 10768 11673 24 NOR2X1 $T=1241540 1465750 1 0 $X=1241538 $Y=1461810
X1710 11744 25 10850 11904 24 NOR2X1 $T=1248900 1480510 0 0 $X=1248898 $Y=1480258
X1711 11904 25 11908 11808 24 NOR2X1 $T=1252120 1473130 1 0 $X=1252118 $Y=1469190
X1712 11937 25 11904 11872 24 NOR2X1 $T=1253960 1473130 1 180 $X=1252580 $Y=1472878
X1713 11948 25 10863 11908 24 NOR2X1 $T=1261320 1473130 0 0 $X=1261318 $Y=1472878
X1714 12075 25 11692 12065 24 NOR2X1 $T=1266840 1487890 1 180 $X=1265460 $Y=1487638
X1715 12183 25 12178 11764 24 NOR2X1 $T=1272360 1473130 0 180 $X=1270980 $Y=1469190
X1716 12065 25 12190 12210 24 NOR2X1 $T=1272360 1473130 0 0 $X=1272358 $Y=1472878
X1717 12222 25 11804 12190 24 NOR2X1 $T=1276500 1480510 0 180 $X=1275120 $Y=1476570
X1718 12315 25 11093 12246 24 NOR2X1 $T=1282020 1465750 1 0 $X=1282018 $Y=1461810
X1719 76 25 10937 12676 24 NOR2X1 $T=1309160 1362430 1 0 $X=1309158 $Y=1358490
X1720 10033 25 10137 12819 24 NOR2X1 $T=1325260 1355050 0 0 $X=1325258 $Y=1354798
X1721 14839 25 386 14921 24 NOR2X1 $T=1526740 1377190 1 0 $X=1526738 $Y=1373250
X1722 512 25 343 547 24 NOR2X1 $T=1528580 1391950 1 180 $X=1527200 $Y=1391698
X1723 14924 25 14874 14844 24 NOR2X1 $T=1530420 1428850 1 180 $X=1529040 $Y=1428598
X1724 14912 25 14870 14856 24 NOR2X1 $T=1530880 1450990 1 180 $X=1529500 $Y=1450738
X1725 374 25 14917 14874 24 NOR2X1 $T=1532720 1436230 1 0 $X=1532718 $Y=1432290
X1726 14924 25 14921 548 24 NOR2X1 $T=1534560 1369810 1 0 $X=1534558 $Y=1365870
X1727 14924 25 14934 14944 24 NOR2X1 $T=1534560 1428850 1 0 $X=1534558 $Y=1424910
X1728 353 25 14833 14945 24 NOR2X1 $T=1535020 1465750 0 0 $X=1535018 $Y=1465498
X1729 547 25 14940 14951 24 NOR2X1 $T=1535480 1391950 0 0 $X=1535478 $Y=1391698
X1730 386 25 14849 14934 24 NOR2X1 $T=1535940 1421470 1 0 $X=1535938 $Y=1417530
X1731 14958 25 14945 14970 24 NOR2X1 $T=1537320 1465750 0 180 $X=1535940 $Y=1461810
X1732 14959 25 14955 14946 24 NOR2X1 $T=1537780 1384570 0 180 $X=1536400 $Y=1380630
X1733 551 25 14956 14931 24 NOR2X1 $T=1537780 1436230 1 180 $X=1536400 $Y=1435978
X1734 15028 25 14950 14954 24 NOR2X1 $T=1538700 1369810 1 180 $X=1537320 $Y=1369558
X1735 549 25 399 551 24 NOR2X1 $T=1537780 1436230 1 0 $X=1537778 $Y=1432290
X1736 551 25 14967 14881 24 NOR2X1 $T=1538240 1428850 1 0 $X=1538238 $Y=1424910
X1737 552 25 357 14912 24 NOR2X1 $T=1538240 1443610 1 0 $X=1538238 $Y=1439670
X1738 554 25 14988 14955 24 NOR2X1 $T=1541460 1384570 0 0 $X=1541458 $Y=1384318
X1739 552 25 383 555 24 NOR2X1 $T=1541920 1428850 0 0 $X=1541918 $Y=1428598
X1740 15051 25 384 14940 24 NOR2X1 $T=1543300 1399330 0 180 $X=1541920 $Y=1395390
X1741 15039 25 554 14967 24 NOR2X1 $T=1543300 1428850 0 180 $X=1541920 $Y=1424910
X1742 14982 25 537 15069 24 NOR2X1 $T=1542380 1495270 0 0 $X=1542378 $Y=1495018
X1743 559 25 14987 14972 24 NOR2X1 $T=1543760 1406710 1 180 $X=1542380 $Y=1406458
X1744 15028 25 15036 14985 24 NOR2X1 $T=1542840 1369810 1 0 $X=1542838 $Y=1365870
X1745 512 25 525 559 24 NOR2X1 $T=1542840 1399330 0 0 $X=1542838 $Y=1399078
X1746 14917 25 554 14956 24 NOR2X1 $T=1542840 1436230 0 0 $X=1542838 $Y=1435978
X1747 512 25 399 14959 24 NOR2X1 $T=1543300 1384570 1 0 $X=1543298 $Y=1380630
X1748 549 25 340 15028 24 NOR2X1 $T=1543300 1458370 1 0 $X=1543298 $Y=1454430
X1749 555 25 15038 14938 24 NOR2X1 $T=1543300 1458370 0 0 $X=1543298 $Y=1458118
X1750 344 25 14982 15038 24 NOR2X1 $T=1543300 1465750 0 0 $X=1543298 $Y=1465498
X1751 14971 25 340 15092 24 NOR2X1 $T=1543300 1473130 1 0 $X=1543298 $Y=1469190
X1752 15030 25 399 15036 24 NOR2X1 $T=1544680 1362430 1 180 $X=1543300 $Y=1362178
X1753 549 25 543 564 24 NOR2X1 $T=1546060 1443610 0 180 $X=1544680 $Y=1439670
X1754 552 25 382 14924 24 NOR2X1 $T=1545140 1428850 0 0 $X=1545138 $Y=1428598
X1755 15028 25 15073 15033 24 NOR2X1 $T=1546520 1465750 1 0 $X=1546518 $Y=1461810
X1756 15127 25 15069 15054 24 NOR2X1 $T=1548360 1495270 1 180 $X=1546980 $Y=1495018
X1757 15030 25 360 15146 24 NOR2X1 $T=1549280 1362430 0 0 $X=1549278 $Y=1362178
X1758 14971 25 344 15147 24 NOR2X1 $T=1549280 1473130 1 0 $X=1549278 $Y=1469190
X1759 569 25 15095 15126 24 NOR2X1 $T=1550660 1369810 1 180 $X=1549280 $Y=1369558
X1760 564 25 15092 15093 24 NOR2X1 $T=1550660 1465750 1 180 $X=1549280 $Y=1465498
X1761 549 25 537 14958 24 NOR2X1 $T=1549740 1450990 0 0 $X=1549738 $Y=1450738
X1762 15028 25 15128 15150 24 NOR2X1 $T=1550200 1450990 1 0 $X=1550198 $Y=1447050
X1763 561 25 15130 15047 24 NOR2X1 $T=1550660 1406710 0 0 $X=1550658 $Y=1406458
X1764 549 25 353 15127 24 NOR2X1 $T=1551120 1495270 0 0 $X=1551118 $Y=1495018
X1765 549 25 343 15140 24 NOR2X1 $T=1551580 1377190 0 0 $X=1551578 $Y=1376938
X1766 552 25 391 561 24 NOR2X1 $T=1552960 1391950 1 0 $X=1552958 $Y=1388010
X1767 15164 25 543 15128 24 NOR2X1 $T=1554800 1443610 0 180 $X=1553420 $Y=1439670
X1768 552 25 386 15158 24 NOR2X1 $T=1554340 1421470 0 0 $X=1554338 $Y=1421218
X1769 570 25 15154 15144 24 NOR2X1 $T=1554340 1502650 1 0 $X=1554338 $Y=1498710
X1770 573 25 15147 15143 24 NOR2X1 $T=1556180 1473130 0 180 $X=1554800 $Y=1469190
X1771 14924 25 15159 15172 24 NOR2X1 $T=1555260 1377190 1 0 $X=1555258 $Y=1373250
X1772 14958 25 15161 15160 24 NOR2X1 $T=1555260 1414090 0 0 $X=1555258 $Y=1413838
X1773 15140 25 15165 15157 24 NOR2X1 $T=1555720 1377190 0 0 $X=1555718 $Y=1376938
X1774 344 25 15166 15168 24 NOR2X1 $T=1555720 1465750 1 0 $X=1555718 $Y=1461810
X1775 15035 25 537 15154 24 NOR2X1 $T=1555720 1495270 0 0 $X=1555718 $Y=1495018
X1776 552 25 374 15170 24 NOR2X1 $T=1556180 1436230 1 0 $X=1556178 $Y=1432290
X1777 549 25 364 570 24 NOR2X1 $T=1556640 1495270 1 0 $X=1556638 $Y=1491330
X1778 15158 25 15146 15156 24 NOR2X1 $T=1557100 1369810 1 0 $X=1557098 $Y=1365870
X1779 15051 25 391 15229 24 NOR2X1 $T=1558940 1391950 0 0 $X=1558938 $Y=1391698
X1780 364 25 15174 15161 24 NOR2X1 $T=1558940 1414090 0 0 $X=1558938 $Y=1413838
X1781 573 25 15184 15190 24 NOR2X1 $T=1558940 1473130 1 0 $X=1558938 $Y=1469190
X1782 15189 25 364 15165 24 NOR2X1 $T=1560320 1377190 1 180 $X=1558940 $Y=1376938
X1783 575 25 386 15226 24 NOR2X1 $T=1560320 1391950 1 0 $X=1560318 $Y=1388010
X1784 15226 25 15229 15193 24 NOR2X1 $T=1561700 1391950 0 0 $X=1561698 $Y=1391698
X1785 552 25 401 580 24 NOR2X1 $T=1561700 1414090 0 0 $X=1561698 $Y=1413838
X1786 15170 25 15232 15285 24 NOR2X1 $T=1562160 1428850 0 0 $X=1562158 $Y=1428598
X1787 580 25 15265 15227 24 NOR2X1 $T=1566760 1436230 0 0 $X=1566758 $Y=1435978
X1788 552 25 360 573 24 NOR2X1 $T=1568140 1428850 1 0 $X=1568138 $Y=1424910
X1789 29 24 25 7872 CLKINVX1 $T=926440 1399330 1 180 $X=925520 $Y=1399078
X1790 31 24 25 9679 CLKINVX1 $T=1079160 1362430 0 180 $X=1078240 $Y=1358490
X1791 34 24 25 9811 CLKINVX1 $T=1092960 1355050 0 0 $X=1092958 $Y=1354798
X1792 45 24 25 9827 CLKINVX1 $T=1097100 1355050 1 180 $X=1096180 $Y=1354798
X1793 9745 24 25 9673 CLKINVX1 $T=1104460 1406710 1 0 $X=1104458 $Y=1402770
X1794 40 24 25 9924 CLKINVX1 $T=1104460 1421470 1 0 $X=1104458 $Y=1417530
X1795 52 24 25 9997 CLKINVX1 $T=1105840 1414090 0 0 $X=1105838 $Y=1413838
X1796 49 24 25 9999 CLKINVX1 $T=1110440 1362430 1 0 $X=1110438 $Y=1358490
X1797 58 24 25 9933 CLKINVX1 $T=1111360 1406710 0 180 $X=1110440 $Y=1402770
X1798 36 24 25 10050 CLKINVX1 $T=1112280 1428850 0 0 $X=1112278 $Y=1428598
X1799 48 24 25 10032 CLKINVX1 $T=1112740 1450990 0 0 $X=1112738 $Y=1450738
X1800 74 24 25 9948 CLKINVX1 $T=1115500 1377190 0 180 $X=1114580 $Y=1373250
X1801 76 24 25 10038 CLKINVX1 $T=1116420 1362430 0 180 $X=1115500 $Y=1358490
X1802 9934 24 25 10117 CLKINVX1 $T=1121940 1421470 0 0 $X=1121938 $Y=1421218
X1803 10004 24 25 10185 CLKINVX1 $T=1127460 1414090 1 0 $X=1127458 $Y=1410150
X1804 10227 24 25 10124 CLKINVX1 $T=1128840 1458370 0 180 $X=1127920 $Y=1454430
X1805 10180 24 25 10186 CLKINVX1 $T=1129300 1458370 1 180 $X=1128380 $Y=1458118
X1806 9995 24 25 10243 CLKINVX1 $T=1129300 1487890 0 0 $X=1129298 $Y=1487638
X1807 9993 24 25 10265 CLKINVX1 $T=1129760 1414090 0 0 $X=1129758 $Y=1413838
X1808 10234 24 25 10143 CLKINVX1 $T=1130680 1465750 1 180 $X=1129760 $Y=1465498
X1809 10261 24 25 10183 CLKINVX1 $T=1130680 1487890 0 180 $X=1129760 $Y=1483950
X1810 10230 24 25 10188 CLKINVX1 $T=1132520 1473130 1 180 $X=1131600 $Y=1472878
X1811 10254 24 25 10238 CLKINVX1 $T=1135280 1458370 1 180 $X=1134360 $Y=1458118
X1812 10266 24 25 10224 CLKINVX1 $T=1136200 1473130 1 180 $X=1135280 $Y=1472878
X1813 10260 24 25 10254 CLKINVX1 $T=1136660 1473130 0 180 $X=1135740 $Y=1469190
X1814 10067 24 25 10273 CLKINVX1 $T=1136200 1414090 1 0 $X=1136198 $Y=1410150
X1815 10263 24 25 10159 CLKINVX1 $T=1138500 1487890 1 0 $X=1138498 $Y=1483950
X1816 10169 24 25 10338 CLKINVX1 $T=1139880 1458370 0 0 $X=1139878 $Y=1458118
X1817 30 24 25 10333 CLKINVX1 $T=1144020 1384570 1 0 $X=1144018 $Y=1380630
X1818 10354 24 25 10287 CLKINVX1 $T=1144940 1436230 1 180 $X=1144020 $Y=1435978
X1819 10359 24 25 10270 CLKINVX1 $T=1145400 1465750 1 180 $X=1144480 $Y=1465498
X1820 10280 24 25 10353 CLKINVX1 $T=1144940 1458370 0 0 $X=1144938 $Y=1458118
X1821 10274 24 25 10386 CLKINVX1 $T=1144940 1487890 1 0 $X=1144938 $Y=1483950
X1822 10343 24 25 10268 CLKINVX1 $T=1146320 1495270 0 180 $X=1145400 $Y=1491330
X1823 10339 24 25 10375 CLKINVX1 $T=1146320 1436230 0 0 $X=1146318 $Y=1435978
X1824 10259 24 25 10483 CLKINVX1 $T=1146780 1465750 1 0 $X=1146778 $Y=1461810
X1825 10226 24 25 10146 CLKINVX1 $T=1148160 1436230 0 180 $X=1147240 $Y=1432290
X1826 10034 24 25 10501 CLKINVX1 $T=1153680 1465750 0 0 $X=1153678 $Y=1465498
X1827 10465 24 25 10473 CLKINVX1 $T=1155520 1487890 0 0 $X=1155518 $Y=1487638
X1828 42 24 25 10587 CLKINVX1 $T=1159200 1428850 0 0 $X=1159198 $Y=1428598
X1829 10594 24 25 10578 CLKINVX1 $T=1161960 1502650 1 180 $X=1161040 $Y=1502398
X1830 120 24 25 10623 CLKINVX1 $T=1161960 1362430 0 0 $X=1161958 $Y=1362178
X1831 10596 24 25 10271 CLKINVX1 $T=1162880 1495270 0 180 $X=1161960 $Y=1491330
X1832 10383 24 25 10607 CLKINVX1 $T=1162880 1377190 1 0 $X=1162878 $Y=1373250
X1833 10360 24 25 10656 CLKINVX1 $T=1162880 1384570 0 0 $X=1162878 $Y=1384318
X1834 10384 24 25 10618 CLKINVX1 $T=1164260 1377190 0 0 $X=1164258 $Y=1376938
X1835 10445 24 25 10619 CLKINVX1 $T=1164260 1391950 1 0 $X=1164258 $Y=1388010
X1836 63 24 25 10632 CLKINVX1 $T=1164260 1436230 0 0 $X=1164258 $Y=1435978
X1837 10480 24 25 10652 CLKINVX1 $T=1167020 1458370 1 0 $X=1167018 $Y=1454430
X1838 10533 24 25 10658 CLKINVX1 $T=1167480 1391950 0 0 $X=1167478 $Y=1391698
X1839 10051 24 25 10676 CLKINVX1 $T=1167480 1465750 0 0 $X=1167478 $Y=1465498
X1840 10464 24 25 10675 CLKINVX1 $T=1168860 1369810 0 0 $X=1168858 $Y=1369558
X1841 10337 24 25 10672 CLKINVX1 $T=1168860 1473130 1 0 $X=1168858 $Y=1469190
X1842 10677 24 25 10712 CLKINVX1 $T=1169780 1465750 1 0 $X=1169778 $Y=1461810
X1843 10535 24 25 10714 CLKINVX1 $T=1170240 1443610 1 0 $X=1170238 $Y=1439670
X1844 10500 24 25 10753 CLKINVX1 $T=1171160 1465750 0 0 $X=1171158 $Y=1465498
X1845 140 24 25 104 CLKINVX1 $T=1172540 1406710 1 180 $X=1171620 $Y=1406458
X1846 119 24 25 10485 CLKINVX1 $T=1173460 1450990 0 0 $X=1173458 $Y=1450738
X1847 132 24 25 10796 CLKINVX1 $T=1173460 1480510 0 0 $X=1173458 $Y=1480258
X1848 10657 24 25 10856 CLKINVX1 $T=1174840 1443610 1 0 $X=1174838 $Y=1439670
X1849 10147 24 25 10774 CLKINVX1 $T=1175300 1465750 0 0 $X=1175298 $Y=1465498
X1850 10814 24 25 10879 CLKINVX1 $T=1179900 1369810 1 0 $X=1179898 $Y=1365870
X1851 10935 24 25 10919 CLKINVX1 $T=1185880 1362430 1 180 $X=1184960 $Y=1362178
X1852 10963 24 25 10971 CLKINVX1 $T=1190020 1369810 0 0 $X=1190018 $Y=1369558
X1853 10711 24 25 11019 CLKINVX1 $T=1190940 1465750 1 0 $X=1190938 $Y=1461810
X1854 10960 24 25 10970 CLKINVX1 $T=1190940 1495270 1 0 $X=1190938 $Y=1491330
X1855 10872 24 25 11027 CLKINVX1 $T=1191860 1377190 0 0 $X=1191858 $Y=1376938
X1856 56 24 25 11023 CLKINVX1 $T=1191860 1458370 1 0 $X=1191858 $Y=1454430
X1857 11015 24 25 10953 CLKINVX1 $T=1192780 1355050 1 180 $X=1191860 $Y=1354798
X1858 69 24 25 11062 CLKINVX1 $T=1192320 1450990 0 0 $X=1192318 $Y=1450738
X1859 10615 24 25 10964 CLKINVX1 $T=1196000 1524790 1 0 $X=1195998 $Y=1520850
X1860 78 24 25 11104 CLKINVX1 $T=1198300 1465750 1 0 $X=1198298 $Y=1461810
X1861 143 24 25 11197 CLKINVX1 $T=1198300 1517410 1 0 $X=1198298 $Y=1513470
X1862 71 24 25 11171 CLKINVX1 $T=1201060 1487890 0 0 $X=1201058 $Y=1487638
X1863 140 24 25 11196 CLKINVX1 $T=1201060 1502650 1 0 $X=1201058 $Y=1498710
X1864 11077 24 25 11107 CLKINVX1 $T=1204740 1355050 1 180 $X=1203820 $Y=1354798
X1865 67 24 25 11213 CLKINVX1 $T=1205200 1458370 0 0 $X=1205198 $Y=1458118
X1866 117 24 25 11223 CLKINVX1 $T=1205200 1502650 1 0 $X=1205198 $Y=1498710
X1867 11117 24 25 11251 CLKINVX1 $T=1207500 1458370 1 0 $X=1207498 $Y=1454430
X1868 64 24 25 11255 CLKINVX1 $T=1209340 1473130 1 0 $X=1209338 $Y=1469190
X1869 11312 24 25 184 CLKINVX1 $T=1210720 1355050 0 180 $X=1209800 $Y=1351110
X1870 11184 24 25 11233 CLKINVX1 $T=1210260 1458370 1 0 $X=1210258 $Y=1454430
X1871 11297 24 25 11357 CLKINVX1 $T=1213480 1369810 1 0 $X=1213478 $Y=1365870
X1872 11368 24 25 10801 CLKINVX1 $T=1219920 1428850 1 180 $X=1219000 $Y=1428598
X1873 11354 24 25 11368 CLKINVX1 $T=1219460 1436230 0 0 $X=1219458 $Y=1435978
X1874 11331 24 25 11388 CLKINVX1 $T=1219920 1377190 1 0 $X=1219918 $Y=1373250
X1875 11073 24 25 11252 CLKINVX1 $T=1221760 1450990 0 0 $X=1221758 $Y=1450738
X1876 195 24 25 11478 CLKINVX1 $T=1222680 1355050 1 0 $X=1222678 $Y=1351110
X1877 11232 24 25 11450 CLKINVX1 $T=1222680 1384570 1 0 $X=1222678 $Y=1380630
X1878 11337 24 25 11489 CLKINVX1 $T=1226360 1369810 0 0 $X=1226358 $Y=1369558
X1879 11520 24 25 11521 CLKINVX1 $T=1228660 1384570 0 0 $X=1228658 $Y=1384318
X1880 11527 24 25 11533 CLKINVX1 $T=1230040 1399330 1 0 $X=1230038 $Y=1395390
X1881 11523 24 25 11580 CLKINVX1 $T=1230500 1458370 1 0 $X=1230498 $Y=1454430
X1882 11477 24 25 11587 CLKINVX1 $T=1230960 1406710 0 0 $X=1230958 $Y=1406458
X1883 11497 24 25 11579 CLKINVX1 $T=1230960 1443610 0 0 $X=1230958 $Y=1443358
X1884 11535 24 25 11618 CLKINVX1 $T=1230960 1473130 1 0 $X=1230958 $Y=1469190
X1885 108 24 25 11596 CLKINVX1 $T=1233720 1502650 1 180 $X=1232800 $Y=1502398
X1886 122 24 25 11585 CLKINVX1 $T=1233260 1495270 1 0 $X=1233258 $Y=1491330
X1887 11543 24 25 11623 CLKINVX1 $T=1234180 1406710 0 0 $X=1234178 $Y=1406458
X1888 11649 24 25 11650 CLKINVX1 $T=1238320 1436230 1 180 $X=1237400 $Y=1435978
X1889 11673 24 25 11743 CLKINVX1 $T=1238780 1465750 1 180 $X=1237860 $Y=1465498
X1890 206 24 25 11600 CLKINVX1 $T=1238320 1355050 0 0 $X=1238318 $Y=1354798
X1891 164 24 25 11179 CLKINVX1 $T=1239700 1443610 1 0 $X=1239698 $Y=1439670
X1892 11678 24 25 11691 CLKINVX1 $T=1242460 1377190 0 180 $X=1241540 $Y=1373250
X1893 11320 24 25 11631 CLKINVX1 $T=1242000 1391950 1 0 $X=1241998 $Y=1388010
X1894 11761 24 25 11620 CLKINVX1 $T=1244300 1532170 1 0 $X=1244298 $Y=1528230
X1895 11773 24 25 221 CLKINVX1 $T=1245220 1355050 1 180 $X=1244300 $Y=1354798
X1896 11899 24 25 234 CLKINVX1 $T=1252120 1362430 0 180 $X=1251200 $Y=1358490
X1897 11904 24 25 11928 CLKINVX1 $T=1254880 1480510 0 0 $X=1254878 $Y=1480258
X1898 11937 24 25 11940 CLKINVX1 $T=1255800 1465750 0 0 $X=1255798 $Y=1465498
X1899 84 24 25 10378 CLKINVX1 $T=1258100 1406710 1 0 $X=1258098 $Y=1402770
X1900 124 24 25 12012 CLKINVX1 $T=1259480 1502650 1 0 $X=1259478 $Y=1498710
X1901 11908 24 25 11933 CLKINVX1 $T=1260860 1465750 0 0 $X=1260858 $Y=1465498
X1902 11897 24 25 11957 CLKINVX1 $T=1263160 1414090 1 0 $X=1263158 $Y=1410150
X1903 12065 24 25 12079 CLKINVX1 $T=1266380 1487890 0 180 $X=1265460 $Y=1483950
X1904 11798 24 25 262 CLKINVX1 $T=1266380 1362430 1 0 $X=1266378 $Y=1358490
X1905 12085 24 25 12181 CLKINVX1 $T=1267300 1421470 0 0 $X=1267298 $Y=1421218
X1906 11877 24 25 263 CLKINVX1 $T=1273280 1362430 0 180 $X=1272360 $Y=1358490
X1907 11252 24 25 11327 CLKINVX1 $T=1277880 1443610 0 0 $X=1277878 $Y=1443358
X1908 11924 24 25 271 CLKINVX1 $T=1278340 1362430 1 0 $X=1278338 $Y=1358490
X1909 12075 24 25 12206 CLKINVX1 $T=1281560 1510030 0 0 $X=1281558 $Y=1509778
X1910 12246 24 25 12262 CLKINVX1 $T=1282480 1458370 0 0 $X=1282478 $Y=1458118
X1911 11662 24 25 12329 CLKINVX1 $T=1282940 1369810 1 0 $X=1282938 $Y=1365870
X1912 11894 24 25 278 CLKINVX1 $T=1283400 1362430 1 0 $X=1283398 $Y=1358490
X1913 11675 24 25 282 CLKINVX1 $T=1283860 1355050 1 0 $X=1283858 $Y=1351110
X1914 11498 24 25 12349 CLKINVX1 $T=1283860 1384570 0 0 $X=1283858 $Y=1384318
X1915 12204 24 25 12055 CLKINVX1 $T=1285240 1406710 1 180 $X=1284320 $Y=1406458
X1916 11792 24 25 291 CLKINVX1 $T=1284780 1377190 1 0 $X=1284778 $Y=1373250
X1917 12313 24 25 287 CLKINVX1 $T=1284780 1384570 1 0 $X=1284778 $Y=1380630
X1918 11617 24 25 276 CLKINVX1 $T=1284780 1458370 0 0 $X=1284778 $Y=1458118
X1919 11620 24 25 12353 CLKINVX1 $T=1285700 1465750 0 180 $X=1284780 $Y=1461810
X1920 12187 24 25 12467 CLKINVX1 $T=1285240 1450990 0 0 $X=1285238 $Y=1450738
X1921 12026 24 25 12384 CLKINVX1 $T=1286620 1428850 0 0 $X=1286618 $Y=1428598
X1922 11463 24 25 12482 CLKINVX1 $T=1290300 1473130 0 0 $X=1290298 $Y=1472878
X1923 11744 24 25 12416 CLKINVX1 $T=1290300 1502650 1 0 $X=1290298 $Y=1498710
X1924 12040 24 25 303 CLKINVX1 $T=1294900 1377190 0 0 $X=1294898 $Y=1376938
X1925 11530 24 25 12490 CLKINVX1 $T=1295360 1421470 1 0 $X=1295358 $Y=1417530
X1926 10391 24 25 12559 CLKINVX1 $T=1296280 1384570 0 0 $X=1296278 $Y=1384318
X1927 11364 24 25 12511 CLKINVX1 $T=1296740 1443610 0 0 $X=1296738 $Y=1443358
X1928 11486 24 25 307 CLKINVX1 $T=1297200 1355050 1 0 $X=1297198 $Y=1351110
X1929 11948 24 25 12565 CLKINVX1 $T=1300420 1517410 1 0 $X=1300418 $Y=1513470
X1930 12500 24 25 12366 CLKINVX1 $T=1301340 1391950 1 0 $X=1301338 $Y=1388010
X1931 12636 24 25 12500 CLKINVX1 $T=1303640 1384570 1 180 $X=1302720 $Y=1384318
X1932 10925 24 25 12608 CLKINVX1 $T=1304560 1391950 0 0 $X=1304558 $Y=1391698
X1933 11496 24 25 12614 CLKINVX1 $T=1305480 1362430 1 0 $X=1305478 $Y=1358490
X1934 10297 24 25 315 CLKINVX1 $T=1308240 1399330 0 0 $X=1308238 $Y=1399078
X1935 12673 24 25 12685 CLKINVX1 $T=1311460 1362430 0 0 $X=1311458 $Y=1362178
X1936 12671 24 25 12793 CLKINVX1 $T=1321120 1369810 1 0 $X=1321118 $Y=1365870
X1937 13294 24 25 304 CLKINVX1 $T=1369880 1473130 1 180 $X=1368960 $Y=1472878
X1938 73 24 25 587 CLKINVX1 $T=1566760 1355050 1 0 $X=1566758 $Y=1351110
X1939 9818 25 24 9828 INVXL $T=1095260 1473130 1 0 $X=1095258 $Y=1469190
X1940 9828 25 24 9934 INVXL $T=1104000 1473130 1 0 $X=1103998 $Y=1469190
X1941 43 25 24 9817 INVXL $T=1105380 1436230 1 180 $X=1104460 $Y=1435978
X1942 9928 25 24 10004 INVXL $T=1105380 1458370 0 0 $X=1105378 $Y=1458118
X1943 9945 25 24 9928 INVXL $T=1106300 1465750 0 180 $X=1105380 $Y=1461810
X1944 9904 25 24 9954 INVXL $T=1109060 1450990 0 0 $X=1109058 $Y=1450738
X1945 60 25 24 9940 INVXL $T=1109980 1384570 0 180 $X=1109060 $Y=1380630
X1946 9954 25 24 10013 INVXL $T=1110900 1450990 0 0 $X=1110898 $Y=1450738
X1947 10007 25 24 10000 INVXL $T=1111820 1465750 1 180 $X=1110900 $Y=1465498
X1948 10052 25 24 9745 INVXL $T=1115960 1436230 0 180 $X=1115040 $Y=1432290
X1949 10000 25 24 10067 INVXL $T=1116420 1465750 0 0 $X=1116418 $Y=1465498
X1950 10073 25 24 10052 INVXL $T=1119180 1436230 0 180 $X=1118260 $Y=1432290
X1951 10155 25 24 10174 INVXL $T=1127460 1473130 0 0 $X=1127458 $Y=1472878
X1952 10173 25 24 90 INVXL $T=1128380 1436230 1 180 $X=1127460 $Y=1435978
X1953 10174 25 24 9993 INVXL $T=1128380 1473130 0 180 $X=1127460 $Y=1469190
X1954 10223 25 24 10173 INVXL $T=1128840 1443610 0 180 $X=1127920 $Y=1439670
X1955 10181 25 24 10169 INVXL $T=1129300 1510030 0 180 $X=1128380 $Y=1506090
X1956 10133 25 24 10181 INVXL $T=1128840 1510030 0 0 $X=1128838 $Y=1509778
X1957 10033 25 24 10249 INVXL $T=1132520 1377190 1 0 $X=1132518 $Y=1373250
X1958 10290 25 24 10180 INVXL $T=1139420 1502650 0 180 $X=1138500 $Y=1498710
X1959 10011 25 24 10290 INVXL $T=1139420 1502650 0 0 $X=1139418 $Y=1502398
X1960 10291 25 24 10299 INVXL $T=1140340 1510030 1 0 $X=1140338 $Y=1506090
X1961 10283 25 24 10370 INVXL $T=1145400 1502650 1 0 $X=1145398 $Y=1498710
X1962 10299 25 24 10369 INVXL $T=1145400 1510030 0 0 $X=1145398 $Y=1509778
X1963 10370 25 24 10280 INVXL $T=1146320 1495270 1 180 $X=1145400 $Y=1495018
X1964 101 25 24 110 INVXL $T=1146780 1355050 1 0 $X=1146778 $Y=1351110
X1965 10388 25 24 10364 INVXL $T=1147700 1414090 0 180 $X=1146780 $Y=1410150
X1966 10503 25 24 10343 INVXL $T=1152300 1510030 1 180 $X=1151380 $Y=1509778
X1967 10491 25 24 10514 INVXL $T=1157360 1502650 1 0 $X=1157358 $Y=1498710
X1968 10470 25 24 10503 INVXL $T=1157360 1510030 0 0 $X=1157358 $Y=1509778
X1969 10514 25 24 10474 INVXL $T=1158280 1495270 1 180 $X=1157360 $Y=1495018
X1970 10589 25 24 10601 INVXL $T=1162420 1406710 1 0 $X=1162418 $Y=1402770
X1971 10588 25 24 10602 INVXL $T=1162420 1421470 1 0 $X=1162418 $Y=1417530
X1972 10591 25 24 10603 INVXL $T=1162420 1421470 0 0 $X=1162418 $Y=1421218
X1973 10600 25 24 10605 INVXL $T=1162880 1502650 0 0 $X=1162878 $Y=1502398
X1974 10511 25 24 10467 INVXL $T=1163800 1480510 1 180 $X=1162880 $Y=1480258
X1975 10610 25 24 10661 INVXL $T=1163800 1399330 1 0 $X=1163798 $Y=1395390
X1976 10581 25 24 10627 INVXL $T=1163800 1510030 0 0 $X=1163798 $Y=1509778
X1977 10648 25 24 10610 INVXL $T=1164720 1399330 1 180 $X=1163800 $Y=1399078
X1978 10605 25 24 10488 INVXL $T=1164720 1502650 0 0 $X=1164718 $Y=1502398
X1979 10627 25 24 10568 INVXL $T=1165180 1510030 1 0 $X=1165178 $Y=1506090
X1980 10601 25 24 10662 INVXL $T=1167480 1406710 1 0 $X=1167478 $Y=1402770
X1981 10602 25 24 10716 INVXL $T=1167480 1421470 1 0 $X=1167478 $Y=1417530
X1982 10603 25 24 10721 INVXL $T=1167480 1421470 0 0 $X=1167478 $Y=1421218
X1983 59 25 24 10391 INVXL $T=1168400 1384570 0 0 $X=1168398 $Y=1384318
X1984 10583 25 24 10373 INVXL $T=1169320 1473130 1 180 $X=1168400 $Y=1472878
X1985 10635 25 24 10708 INVXL $T=1169320 1428850 0 0 $X=1169318 $Y=1428598
X1986 10708 25 24 10794 INVXL $T=1174380 1428850 0 0 $X=1174378 $Y=1428598
X1987 10763 25 24 10812 INVXL $T=1178980 1510030 0 0 $X=1178978 $Y=1509778
X1988 10629 25 24 10862 INVXL $T=1179900 1458370 1 0 $X=1179898 $Y=1454430
X1989 10671 25 24 10877 INVXL $T=1181280 1443610 1 0 $X=1181278 $Y=1439670
X1990 10877 25 24 10897 INVXL $T=1182200 1436230 0 0 $X=1182198 $Y=1435978
X1991 10812 25 24 10882 INVXL $T=1182660 1510030 0 0 $X=1182658 $Y=1509778
X1992 10911 25 24 10923 INVXL $T=1184040 1480510 0 0 $X=1184038 $Y=1480258
X1993 10923 25 24 10892 INVXL $T=1185880 1487890 1 0 $X=1185878 $Y=1483950
X1994 156 25 24 10930 INVXL $T=1186800 1369810 0 180 $X=1185880 $Y=1365870
X1995 10861 25 24 11016 INVXL $T=1186340 1377190 0 0 $X=1186338 $Y=1376938
X1996 10894 25 24 11030 INVXL $T=1191860 1473130 1 0 $X=1191858 $Y=1469190
X1997 10802 25 24 11056 INVXL $T=1196460 1458370 0 0 $X=1196458 $Y=1458118
X1998 10938 25 24 11064 INVXL $T=1196920 1414090 0 0 $X=1196918 $Y=1413838
X1999 11030 25 24 11163 INVXL $T=1196920 1473130 1 0 $X=1196918 $Y=1469190
X2000 11064 25 24 11188 INVXL $T=1198300 1406710 1 0 $X=1198298 $Y=1402770
X2001 11082 25 24 11100 INVXL $T=1198300 1406710 0 0 $X=1198298 $Y=1406458
X2002 11056 25 24 11075 INVXL $T=1198300 1450990 1 0 $X=1198298 $Y=1447050
X2003 11100 25 24 11079 INVXL $T=1200600 1406710 0 0 $X=1200598 $Y=1406458
X2004 11071 25 24 11323 INVXL $T=1205660 1532170 1 0 $X=1205658 $Y=1528230
X2005 11260 25 24 11253 INVXL $T=1210720 1480510 1 180 $X=1209800 $Y=1480258
X2006 11235 25 24 11306 INVXL $T=1212100 1502650 1 0 $X=1212098 $Y=1498710
X2007 11253 25 24 11308 INVXL $T=1212560 1480510 0 0 $X=1212558 $Y=1480258
X2008 11126 25 24 11329 INVXL $T=1213480 1414090 1 0 $X=1213478 $Y=1410150
X2009 11060 25 24 11355 INVXL $T=1213480 1495270 1 0 $X=1213478 $Y=1491330
X2010 11346 25 24 11334 INVXL $T=1215780 1532170 0 180 $X=1214860 $Y=1528230
X2011 11329 25 24 11393 INVXL $T=1215320 1414090 0 0 $X=1215318 $Y=1413838
X2012 11306 25 24 11364 INVXL $T=1217160 1502650 1 0 $X=1217158 $Y=1498710
X2013 11314 25 24 11397 INVXL $T=1219000 1421470 0 0 $X=1218998 $Y=1421218
X2014 11339 25 24 11475 INVXL $T=1220380 1391950 1 0 $X=1220378 $Y=1388010
X2015 111 25 24 11222 INVXL $T=1221760 1517410 1 0 $X=1221758 $Y=1513470
X2016 11355 25 24 11430 INVXL $T=1222680 1495270 1 0 $X=1222678 $Y=1491330
X2017 11334 25 24 11463 INVXL $T=1223600 1532170 1 0 $X=1223598 $Y=1528230
X2018 11482 25 24 11477 INVXL $T=1225900 1406710 1 180 $X=1224980 $Y=1406458
X2019 11323 25 24 11369 INVXL $T=1225440 1524790 0 0 $X=1225438 $Y=1524538
X2020 11397 25 24 11583 INVXL $T=1232800 1421470 0 0 $X=1232798 $Y=1421218
X2021 11582 25 24 11659 INVXL $T=1237400 1399330 0 0 $X=1237398 $Y=1399078
X2022 11502 25 24 11735 INVXL $T=1237860 1436230 1 0 $X=1237858 $Y=1432290
X2023 11539 25 24 11761 INVXL $T=1241540 1532170 0 0 $X=1241538 $Y=1531918
X2024 100 25 24 11685 INVXL $T=1242460 1502650 1 0 $X=1242458 $Y=1498710
X2025 11769 25 24 11736 INVXL $T=1243380 1414090 0 180 $X=1242460 $Y=1410150
X2026 11588 25 24 11697 INVXL $T=1242920 1362430 1 0 $X=1242918 $Y=1358490
X2027 11784 25 24 11499 INVXL $T=1243840 1458370 0 180 $X=1242920 $Y=1454430
X2028 11624 25 24 11769 INVXL $T=1244300 1414090 0 0 $X=1244298 $Y=1413838
X2029 11653 25 24 11741 INVXL $T=1244760 1377190 1 0 $X=1244758 $Y=1373250
X2030 95 25 24 11888 INVXL $T=1247980 1495270 1 0 $X=1247978 $Y=1491330
X2031 11811 25 24 11801 INVXL $T=1248900 1436230 1 180 $X=1247980 $Y=1435978
X2032 11772 25 24 11870 INVXL $T=1248900 1532170 0 0 $X=1248898 $Y=1531918
X2033 11805 25 24 11812 INVXL $T=1249820 1480510 0 180 $X=1248900 $Y=1476570
X2034 11870 25 24 11744 INVXL $T=1249820 1524790 0 180 $X=1248900 $Y=1520850
X2035 88 25 24 11886 INVXL $T=1250280 1502650 0 0 $X=1250278 $Y=1502398
X2036 11803 25 24 11906 INVXL $T=1251200 1532170 1 0 $X=1251198 $Y=1528230
X2037 11906 25 24 11948 INVXL $T=1254420 1524790 1 0 $X=1254418 $Y=1520850
X2038 11941 25 24 235 INVXL $T=1256720 1406710 1 180 $X=1255800 $Y=1406458
X2039 11764 25 24 11885 INVXL $T=1257180 1473130 0 180 $X=1256260 $Y=1469190
X2040 12033 25 24 11941 INVXL $T=1261780 1406710 1 180 $X=1260860 $Y=1406458
X2041 11801 25 24 12026 INVXL $T=1261320 1436230 0 0 $X=1261318 $Y=1435978
X2042 11895 25 24 12039 INVXL $T=1261780 1539550 1 0 $X=1261778 $Y=1535610
X2043 65 25 24 12062 INVXL $T=1264540 1502650 1 0 $X=1264538 $Y=1498710
X2044 12078 25 24 12016 INVXL $T=1265920 1428850 0 180 $X=1265000 $Y=1424910
X2045 12036 25 24 12076 INVXL $T=1265920 1443610 1 0 $X=1265918 $Y=1439670
X2046 12034 25 24 11784 INVXL $T=1266380 1443610 0 0 $X=1266378 $Y=1443358
X2047 12060 25 24 12078 INVXL $T=1267300 1428850 1 0 $X=1267298 $Y=1424910
X2048 12039 25 24 12075 INVXL $T=1268220 1539550 1 0 $X=1268218 $Y=1535610
X2049 12076 25 24 12187 INVXL $T=1270980 1443610 1 0 $X=1270978 $Y=1439670
X2050 11784 25 24 12189 INVXL $T=1272360 1443610 0 0 $X=1272358 $Y=1443358
X2051 12217 25 24 12185 INVXL $T=1275120 1465750 0 180 $X=1274200 $Y=1461810
X2052 12037 25 24 12234 INVXL $T=1276960 1539550 1 0 $X=1276958 $Y=1535610
X2053 12190 25 24 12242 INVXL $T=1278340 1473130 0 0 $X=1278338 $Y=1472878
X2054 12229 25 24 12247 INVXL $T=1278800 1517410 0 0 $X=1278798 $Y=1517158
X2055 12234 25 24 12222 INVXL $T=1278800 1532170 0 0 $X=1278798 $Y=1531918
X2056 12327 25 24 12335 INVXL $T=1282480 1421470 0 0 $X=1282478 $Y=1421218
X2057 12322 25 24 12338 INVXL $T=1282940 1524790 0 0 $X=1282938 $Y=1524538
X2058 12338 25 24 12201 INVXL $T=1283400 1524790 1 0 $X=1283398 $Y=1520850
X2059 12343 25 24 12352 INVXL $T=1283860 1532170 0 0 $X=1283858 $Y=1531918
X2060 12335 25 24 11662 INVXL $T=1284780 1421470 0 0 $X=1284778 $Y=1421218
X2061 12314 25 24 12367 INVXL $T=1285240 1414090 0 0 $X=1285238 $Y=1413838
X2062 12367 25 24 220 INVXL $T=1286160 1399330 1 180 $X=1285240 $Y=1399078
X2063 12352 25 24 12315 INVXL $T=1288920 1532170 0 0 $X=1288918 $Y=1531918
X2064 12208 25 24 12414 INVXL $T=1290300 1406710 0 0 $X=1290298 $Y=1406458
X2065 12201 25 24 12415 INVXL $T=1290300 1487890 0 0 $X=1290298 $Y=1487638
X2066 12222 25 24 12505 INVXL $T=1295360 1517410 0 0 $X=1295358 $Y=1517158
X2067 12414 25 24 11498 INVXL $T=1296280 1406710 0 0 $X=1296278 $Y=1406458
X2068 12315 25 24 12584 INVXL $T=1302720 1495270 1 0 $X=1302718 $Y=1491330
X2069 68 25 24 12812 INVXL $T=1328480 1362430 0 0 $X=1328478 $Y=1362178
X2070 14839 25 24 14852 INVXL $T=1524900 1362430 1 0 $X=1524898 $Y=1358490
X2071 14833 25 24 14858 INVXL $T=1526740 1480510 0 0 $X=1526738 $Y=1480258
X2072 14849 25 24 14929 INVXL $T=1527200 1421470 1 0 $X=1527198 $Y=1417530
X2073 15035 25 24 14986 INVXL $T=1542380 1495270 0 180 $X=1541460 $Y=1491330
X2074 15039 25 24 15068 INVXL $T=1547900 1406710 1 180 $X=1546980 $Y=1406458
X2075 15164 25 24 15090 INVXL $T=1556640 1436230 1 180 $X=1555720 $Y=1435978
X2076 15174 25 24 15138 INVXL $T=1559860 1421470 0 0 $X=1559858 $Y=1421218
X2077 15166 25 24 15240 INVXL $T=1559860 1480510 0 0 $X=1559858 $Y=1480258
X2078 14988 25 24 15244 INVXL $T=1562620 1384570 0 0 $X=1562618 $Y=1384318
X2079 9926 24 25 9908 INVX1 $T=1104920 1362430 0 180 $X=1104000 $Y=1358490
X2080 10364 24 25 105 INVX1 $T=1141720 1391950 1 180 $X=1140800 $Y=1391698
X2081 10371 24 25 10267 INVX1 $T=1148620 1480510 0 0 $X=1148618 $Y=1480258
X2082 10505 24 25 10389 INVX1 $T=1159200 1473130 0 180 $X=1158280 $Y=1469190
X2083 10614 24 25 10492 INVX1 $T=1169320 1480510 1 180 $X=1168400 $Y=1480258
X2084 151 24 25 10772 INVX1 $T=1180820 1355050 1 180 $X=1179900 $Y=1354798
X2085 10817 24 25 11220 INVX1 $T=1203820 1450990 0 0 $X=1203818 $Y=1450738
X2086 186 24 25 11336 INVX1 $T=1208880 1355050 0 0 $X=1208878 $Y=1354798
X2087 11215 24 25 11262 INVX1 $T=1210720 1510030 1 0 $X=1210718 $Y=1506090
X2088 11123 24 25 11105 INVX1 $T=1214860 1480510 0 0 $X=1214858 $Y=1480258
X2089 11350 24 25 11469 INVX1 $T=1216240 1406710 0 0 $X=1216238 $Y=1406458
X2090 11509 24 25 11452 INVX1 $T=1228200 1428850 1 180 $X=1227280 $Y=1428598
X2091 11441 24 25 11543 INVX1 $T=1232800 1428850 0 0 $X=1232798 $Y=1428598
X2092 11754 24 25 11588 INVX1 $T=1243840 1355050 1 180 $X=1242920 $Y=1354798
X2093 11763 24 25 11770 INVX1 $T=1244300 1443610 1 0 $X=1244298 $Y=1439670
X2094 11871 24 25 11800 INVX1 $T=1249820 1391950 0 180 $X=1248900 $Y=1388010
X2095 11932 24 25 11881 INVX1 $T=1252580 1436230 1 180 $X=1251660 $Y=1435978
X2096 11873 24 25 11958 INVX1 $T=1257640 1421470 0 0 $X=1257638 $Y=1421218
X2097 12168 24 25 12061 INVX1 $T=1267300 1450990 1 180 $X=1266380 $Y=1450738
X2098 12179 24 25 12073 INVX1 $T=1270520 1487890 0 180 $X=1269600 $Y=1483950
X2099 12254 24 25 12333 INVX1 $T=1280180 1436230 1 0 $X=1280178 $Y=1432290
X2100 12243 24 25 12017 INVX1 $T=1282940 1495270 1 0 $X=1282938 $Y=1491330
X2101 101 24 25 10937 INVX1 $T=1285240 1458370 1 0 $X=1285238 $Y=1454430
X2102 543 24 25 14851 INVX1 $T=1525820 1369810 0 0 $X=1525818 $Y=1369558
X2103 340 24 25 15041 INVX1 $T=1544680 1473130 0 0 $X=1544678 $Y=1472878
X2104 357 24 25 15142 INVX1 $T=1552960 1428850 0 0 $X=1552958 $Y=1428598
X2105 15152 24 25 15162 INVX1 $T=1555260 1458370 1 0 $X=1555258 $Y=1454430
X2106 386 24 25 15191 INVX1 $T=1559860 1443610 1 0 $X=1559858 $Y=1439670
X2107 391 24 25 15183 INVX1 $T=1560780 1473130 1 180 $X=1559860 $Y=1472878
X2108 9907 24 10297 25 CLKINVX3 $T=1138040 1414090 0 0 $X=1138038 $Y=1413838
X2109 10126 24 157 25 CLKINVX3 $T=1174840 1391950 0 0 $X=1174838 $Y=1391698
X2110 11626 24 285 25 CLKINVX3 $T=1277880 1450990 0 0 $X=1277878 $Y=1450738
X2111 11917 24 297 25 CLKINVX3 $T=1287540 1355050 0 0 $X=1287538 $Y=1354798
X2112 304 24 11487 25 CLKINVX3 $T=1295360 1473130 0 0 $X=1295358 $Y=1472878
X2113 575 24 562 25 CLKINVX3 $T=1556640 1399330 1 180 $X=1555260 $Y=1399078
X2114 24 25 568 ANTENNA $T=1550660 1546930 1 0 $X=1550658 $Y=1542990
X2115 328 24 10298 25 CLKBUFX20 $T=1328940 1406710 1 0 $X=1328938 $Y=1402770
X2116 328 24 14144 25 CLKBUFX20 $T=1548820 1642870 1 0 $X=1548818 $Y=1638930
X2117 25 12489 308 12561 12388 24 12370 12593 12619 11960 322 12497 12526 12707 3961 ICV_28 $T=1301800 1539550 0 0 $X=1301798 $Y=1539298
X2118 25 12525 300 12595 12582 24 11874 12617 12595 12113 322 12560 12582 12694 3961 ICV_28 $T=1302260 1458370 0 0 $X=1302258 $Y=1458118
X2119 25 12528 299 12609 12602 24 12478 12621 12625 12113 322 12687 12672 12701 3961 ICV_28 $T=1302720 1414090 0 0 $X=1302718 $Y=1413838
X2120 25 12525 305 12598 12403 24 12054 12463 12623 12113 327 12615 12590 12717 3961 ICV_28 $T=1302720 1480510 1 0 $X=1302718 $Y=1476570
X2121 25 12489 299 12622 12621 24 12478 12627 12622 12113 327 12398 12621 12725 3961 ICV_28 $T=1304560 1428850 1 0 $X=1304558 $Y=1424910
X2122 25 12528 311 12779 12782 24 289 12780 12779 229 325 12507 12782 12875 3961 ICV_28 $T=1318820 1391950 1 0 $X=1318818 $Y=1388010
X2123 25 12489 313 12691 12715 24 12370 12801 12809 11960 12641 12721 12896 12969 3961 ICV_28 $T=1319740 1524790 1 0 $X=1319738 $Y=1520850
X2124 25 12806 299 12823 12829 24 12478 12836 12823 229 348 12462 12829 12958 3961 ICV_28 $T=1324800 1414090 1 0 $X=1324798 $Y=1410150
X2125 25 13313 300 13438 13395 24 13294 13395 13486 13102 13225 13576 13533 13584 3961 ICV_28 $T=1379540 1465750 1 0 $X=1379538 $Y=1461810
X2126 25 13313 310 13480 13484 24 12942 13477 13480 13102 13225 12926 13484 13586 3961 ICV_28 $T=1380920 1399330 0 0 $X=1380918 $Y=1399078
X2127 25 461 299 13710 13714 24 13704 13714 13674 13102 454 13383 13689 13823 3961 ICV_28 $T=1405760 1428850 0 0 $X=1405758 $Y=1428598
X2128 25 464 301 13845 13848 24 13789 13864 13845 13368 457 13062 13848 13762 3961 ICV_28 $T=1421400 1532170 0 0 $X=1421398 $Y=1531918
X2129 25 461 312 13856 13847 24 13704 13847 13879 13766 475 12508 13851 13958 3961 ICV_28 $T=1423240 1450990 1 0 $X=1423238 $Y=1447050
X2130 25 13826 313 14241 14243 24 14194 14252 14241 14256 469 13042 14243 14415 3961 ICV_28 $T=1459120 1524790 0 0 $X=1459118 $Y=1524538
X2131 25 13885 14356 14470 14468 24 14282 14554 14559 14370 502 13503 14649 14540 3961 ICV_28 $T=1491780 1421470 1 0 $X=1491778 $Y=1417530
X2132 25 14318 14467 14680 14684 24 14446 14693 14680 14256 14228 13096 14684 14786 3961 ICV_28 $T=1506500 1517410 1 0 $X=1506498 $Y=1513470
X2133 25 14318 14255 14872 14873 24 14446 14837 14872 14256 14228 13096 14873 14832 3961 ICV_28 $T=1526740 1510030 0 0 $X=1526738 $Y=1509778
X2134 25 14859 13891 15043 15060 24 14659 15064 15043 530 453 13476 15060 14988 3961 ICV_28 $T=1542840 1384570 0 0 $X=1542838 $Y=1384318
X2135 12694 12711 334 12385 12740 339 24 12797 25 MXI4X1 $T=1315140 1465750 1 0 $X=1315138 $Y=1461810
X2136 12695 12712 12718 12728 12741 340 24 12798 25 MXI4X1 $T=1315140 1495270 1 0 $X=1315138 $Y=1491330
X2137 12701 12680 12724 12410 12739 342 24 12807 25 MXI4X1 $T=1316060 1399330 0 0 $X=1316058 $Y=1399078
X2138 12634 12725 12729 12383 12706 12802 24 12814 25 MXI4X1 $T=1316520 1421470 1 0 $X=1316518 $Y=1417530
X2139 12708 12516 12733 12732 12677 12811 24 12813 25 MXI4X1 $T=1316980 1532170 1 0 $X=1316978 $Y=1528230
X2140 12703 12730 12734 12520 12698 343 24 12816 25 MXI4X1 $T=1316980 1539550 0 0 $X=1316978 $Y=1539298
X2141 12703 12730 12735 12520 12698 12811 24 12893 25 MXI4X1 $T=1316980 1546930 0 0 $X=1316978 $Y=1546678
X2142 12694 12711 335 12385 12740 344 24 12817 25 MXI4X1 $T=1317440 1458370 0 0 $X=1317438 $Y=1458118
X2143 12690 12717 12718 12626 12783 12802 24 12837 25 MXI4X1 $T=1319280 1487890 0 0 $X=1319278 $Y=1487638
X2144 12707 12669 12735 12331 12786 12811 24 12899 25 MXI4X1 $T=1319280 1539550 1 0 $X=1319278 $Y=1535610
X2145 12690 12717 12788 12626 12783 347 24 12891 25 MXI4X1 $T=1319740 1480510 0 0 $X=1319738 $Y=1480258
X2146 12701 12680 12790 12410 12739 12828 24 12832 25 MXI4X1 $T=1320200 1406710 1 0 $X=1320198 $Y=1402770
X2147 12710 12731 12729 12594 12745 12802 24 12882 25 MXI4X1 $T=1320200 1450990 1 0 $X=1320198 $Y=1447050
X2148 12695 12712 12788 12728 12741 12811 24 12880 25 MXI4X1 $T=1321580 1502650 1 0 $X=1321578 $Y=1498710
X2149 12708 12516 12810 12732 12677 353 24 12892 25 MXI4X1 $T=1322040 1524790 0 0 $X=1322038 $Y=1524538
X2150 12742 12808 12810 12784 12791 12802 24 12845 25 MXI4X1 $T=1322500 1502650 0 0 $X=1322498 $Y=1502398
X2151 12710 12731 12820 12594 12745 344 24 12918 25 MXI4X1 $T=1323880 1443610 0 0 $X=1323878 $Y=1443358
X2152 12772 12689 345 12569 12697 356 24 12890 25 MXI4X1 $T=1323880 1450990 0 0 $X=1323878 $Y=1450738
X2153 12742 12808 12733 12784 12791 356 24 12923 25 MXI4X1 $T=1323880 1510030 1 0 $X=1323878 $Y=1506090
X2154 12723 12824 12820 12521 12719 358 24 12887 25 MXI4X1 $T=1325260 1369810 0 0 $X=1325258 $Y=1369558
X2155 12634 12725 12820 12383 12706 360 24 12922 25 MXI4X1 $T=1325260 1421470 1 0 $X=1325258 $Y=1417530
X2156 12707 12669 12734 12331 12786 353 24 12900 25 MXI4X1 $T=1325720 1539550 0 0 $X=1325718 $Y=1539298
X2157 12772 12689 351 12569 12697 364 24 12903 25 MXI4X1 $T=1326180 1458370 0 0 $X=1326178 $Y=1458118
X2158 12821 12834 352 12714 12875 357 24 12905 25 MXI4X1 $T=1326640 1384570 0 0 $X=1326638 $Y=1384318
X2159 12723 12824 12729 12521 12719 367 24 13033 25 MXI4X1 $T=1327100 1377190 1 0 $X=1327098 $Y=1373250
X2160 349 350 354 319 361 367 24 12915 25 MXI4X1 $T=1328020 1355050 1 0 $X=1328018 $Y=1351110
X2161 12838 12704 12790 12727 12889 12828 24 12932 25 MXI4X1 $T=1328940 1421470 0 0 $X=1328938 $Y=1421218
X2162 12838 12704 12724 12727 12889 342 24 12971 25 MXI4X1 $T=1329860 1428850 0 0 $X=1329858 $Y=1428598
X2163 12821 12834 359 12714 12875 373 24 12959 25 MXI4X1 $T=1330320 1384570 1 0 $X=1330318 $Y=1380630
X2164 12902 12908 12790 12943 12966 12828 24 12970 25 MXI4X1 $T=1335380 1428850 1 0 $X=1335378 $Y=1424910
X2165 12885 12913 345 12950 12964 356 24 13021 25 MXI4X1 $T=1335380 1465750 0 0 $X=1335378 $Y=1465498
X2166 12878 12952 12733 12969 12815 356 24 13031 25 MXI4X1 $T=1337220 1517410 0 0 $X=1337218 $Y=1517158
X2167 12902 12908 12724 12943 12966 342 24 13058 25 MXI4X1 $T=1340900 1428850 0 0 $X=1340898 $Y=1428598
X2168 12885 12913 351 12950 12964 384 24 13111 25 MXI4X1 $T=1340900 1473130 1 0 $X=1340898 $Y=1469190
X2169 12878 12952 12810 12969 12815 373 24 13059 25 MXI4X1 $T=1340900 1517410 1 0 $X=1340898 $Y=1513470
X2170 12792 12946 12735 13026 13037 12811 24 13063 25 MXI4X1 $T=1340900 1539550 0 0 $X=1340898 $Y=1539298
X2171 12792 12946 12734 13026 13037 340 24 13098 25 MXI4X1 $T=1342740 1546930 1 0 $X=1342738 $Y=1542990
X2172 12975 13036 12788 13024 13022 12811 24 13100 25 MXI4X1 $T=1344120 1502650 0 0 $X=1344118 $Y=1502398
X2173 12975 13036 12718 13024 13022 373 24 13116 25 MXI4X1 $T=1344580 1495270 0 0 $X=1344578 $Y=1495018
X2174 12912 12577 12790 13105 13046 365 24 13151 25 MXI4X1 $T=1348260 1399330 0 0 $X=1348258 $Y=1399078
X2175 12912 12577 12724 13105 13046 342 24 13161 25 MXI4X1 $T=1349180 1406710 1 0 $X=1349178 $Y=1402770
X2176 13158 13140 12820 13120 12958 386 24 13054 25 MXI4X1 $T=1357920 1414090 0 180 $X=1349180 $Y=1410150
X2177 12833 13133 12733 13050 13034 356 24 13060 25 MXI4X1 $T=1357920 1524790 1 180 $X=1349180 $Y=1524538
X2178 387 388 354 392 395 367 24 13175 25 MXI4X1 $T=1351020 1355050 1 0 $X=1351018 $Y=1351110
X2179 12939 13016 12820 13094 13147 398 24 13176 25 MXI4X1 $T=1351020 1369810 0 0 $X=1351018 $Y=1369558
X2180 13032 13103 345 13131 13106 12828 24 13178 25 MXI4X1 $T=1351020 1450990 0 0 $X=1351018 $Y=1450738
X2181 13066 12944 12718 13132 12973 12802 24 13171 25 MXI4X1 $T=1351020 1495270 1 0 $X=1351018 $Y=1491330
X2182 13165 13159 12733 13145 13129 356 24 13097 25 MXI4X1 $T=1359760 1539550 0 180 $X=1351020 $Y=1535610
X2183 13099 13118 12734 13110 13017 399 24 13183 25 MXI4X1 $T=1351480 1546930 1 0 $X=1351478 $Y=1542990
X2184 13099 13118 12735 13110 13017 12811 24 13169 25 MXI4X1 $T=1351480 1546930 0 0 $X=1351478 $Y=1546678
X2185 13032 13103 351 13131 13106 342 24 13185 25 MXI4X1 $T=1351940 1458370 1 0 $X=1351938 $Y=1454430
X2186 13109 13119 359 13049 13028 373 24 13189 25 MXI4X1 $T=1352400 1384570 0 0 $X=1352398 $Y=1384318
X2187 12939 13016 12729 13094 13147 367 24 13216 25 MXI4X1 $T=1352860 1377190 1 0 $X=1352858 $Y=1373250
X2188 13114 13124 12788 13095 13113 357 24 13217 25 MXI4X1 $T=1352860 1443610 0 0 $X=1352858 $Y=1443358
X2189 13066 12944 12788 13132 12973 401 24 13168 25 MXI4X1 $T=1352860 1480510 0 0 $X=1352858 $Y=1480258
X2190 12833 13133 12810 13050 13034 12802 24 13218 25 MXI4X1 $T=1352860 1532170 1 0 $X=1352858 $Y=1528230
X2191 13158 13140 12729 13120 12958 12802 24 13130 25 MXI4X1 $T=1363440 1414090 1 180 $X=1354700 $Y=1413838
X2192 13114 13124 12718 13095 13113 12802 24 13273 25 MXI4X1 $T=1355160 1450990 1 0 $X=1355158 $Y=1447050
X2193 13109 13119 352 13049 13028 386 24 13268 25 MXI4X1 $T=1358380 1391950 1 0 $X=1358378 $Y=1388010
X2194 13289 13264 30 12887 13176 396 24 13184 25 MXI4X1 $T=1368500 1369810 1 180 $X=1359760 $Y=1369558
X2195 13308 13282 12724 13260 13244 342 24 13162 25 MXI4X1 $T=1369880 1428850 0 180 $X=1361140 $Y=1424910
X2196 13308 13282 12790 13260 13244 12828 24 13038 25 MXI4X1 $T=1370340 1421470 1 180 $X=1361600 $Y=1421218
X2197 13401 13378 12734 13353 13309 384 24 13172 25 MXI4X1 $T=1375860 1502650 1 180 $X=1367120 $Y=1502398
X2198 13402 13379 12735 13317 13310 12811 24 13135 25 MXI4X1 $T=1375860 1539550 1 180 $X=1367120 $Y=1539298
X2199 13405 13384 12718 13359 13316 12802 24 13246 25 MXI4X1 $T=1376320 1487890 1 180 $X=1367580 $Y=1487638
X2200 13315 13396 351 13373 13351 399 24 13235 25 MXI4X1 $T=1377240 1473130 0 180 $X=1368500 $Y=1469190
X2201 13402 13379 12734 13317 13310 340 24 13262 25 MXI4X1 $T=1377700 1546930 0 180 $X=1368960 $Y=1542990
X2202 13416 13407 433 12832 13151 418 24 13297 25 MXI4X1 $T=1378620 1399330 1 180 $X=1369880 $Y=1399078
X2203 13315 13396 345 13373 13351 356 24 13163 25 MXI4X1 $T=1378620 1465750 0 180 $X=1369880 $Y=1461810
X2204 13401 13378 12735 13353 13309 12811 24 13164 25 MXI4X1 $T=1378620 1510030 0 180 $X=1369880 $Y=1506090
X2205 13398 13375 12733 13322 13305 356 24 13277 25 MXI4X1 $T=1379540 1517410 0 180 $X=1370800 $Y=1513470
X2206 13405 13384 12788 13359 13316 401 24 13236 25 MXI4X1 $T=1380460 1487890 0 180 $X=1371720 $Y=1483950
X2207 13490 13427 12729 13417 13410 12802 24 13255 25 MXI4X1 $T=1382300 1414090 1 180 $X=1373560 $Y=1413838
X2208 13443 13432 12820 13318 13415 398 24 13289 25 MXI4X1 $T=1383220 1369810 1 180 $X=1374480 $Y=1369558
X2209 13482 13433 12718 13424 13370 12802 24 13392 25 MXI4X1 $T=1383220 1443610 1 180 $X=1374480 $Y=1443358
X2210 13443 13432 12729 13318 13415 367 24 13274 25 MXI4X1 $T=1384140 1377190 0 180 $X=1375400 $Y=1373250
X2211 13490 13427 12820 13417 13410 360 24 13148 25 MXI4X1 $T=1384140 1421470 1 180 $X=1375400 $Y=1421218
X2212 13482 13433 12788 13424 13370 374 24 13275 25 MXI4X1 $T=1384600 1443610 0 180 $X=1375860 $Y=1439670
X2213 13497 13487 13143 12900 13183 400 24 13352 25 MXI4X1 $T=1386440 1546930 0 180 $X=1377700 $Y=1542990
X2214 13524 13471 442 13473 13489 391 24 13404 25 MXI4X1 $T=1390120 1391950 0 180 $X=1381380 $Y=1388010
X2215 13524 13471 444 13473 13489 384 24 13271 25 MXI4X1 $T=1390580 1384570 1 180 $X=1381840 $Y=1384318
X2216 449 445 354 443 440 367 24 13293 25 MXI4X1 $T=1391960 1355050 0 180 $X=1383220 $Y=1351110
X2217 13505 13511 12735 13520 13507 12811 24 13239 25 MXI4X1 $T=1392880 1546930 1 180 $X=1384140 $Y=1546678
X2218 13505 13511 12734 13520 13507 384 24 13497 25 MXI4X1 $T=1395180 1546930 0 180 $X=1386440 $Y=1542990
X2219 13657 13589 12718 13577 13535 12802 24 13224 25 MXI4X1 $T=1397020 1487890 1 180 $X=1388280 $Y=1487638
X2220 13624 13613 12790 13488 13586 365 24 13416 25 MXI4X1 $T=1400240 1399330 0 180 $X=1391500 $Y=1395390
X2221 13527 13588 345 13595 13584 12828 24 13256 25 MXI4X1 $T=1392880 1450990 0 0 $X=1392878 $Y=1450738
X2222 13527 13588 351 13595 13584 342 24 13393 25 MXI4X1 $T=1392880 1458370 0 0 $X=1392878 $Y=1458118
X2223 13662 13528 345 13608 13600 356 24 13142 25 MXI4X1 $T=1401620 1465750 1 180 $X=1392880 $Y=1465498
X2224 13657 13589 12788 13577 13535 382 24 13220 25 MXI4X1 $T=1401620 1487890 0 180 $X=1392880 $Y=1483950
X2225 13664 13623 12810 13609 13602 373 24 13221 25 MXI4X1 $T=1401620 1510030 1 180 $X=1392880 $Y=1509778
X2226 13665 13627 12820 13617 13604 358 24 13264 25 MXI4X1 $T=1402540 1369810 1 180 $X=1393800 $Y=1369558
X2227 13670 13652 12734 13626 13618 343 24 13487 25 MXI4X1 $T=1403920 1546930 0 180 $X=1395180 $Y=1542990
X2228 13522 13614 12729 13625 13656 12802 24 13372 25 MXI4X1 $T=1396100 1443610 0 0 $X=1396098 $Y=1443358
X2229 13624 13613 12724 13488 13586 342 24 13243 25 MXI4X1 $T=1404840 1399330 1 180 $X=1396100 $Y=1399078
X2230 13662 13528 351 13608 13600 353 24 13219 25 MXI4X1 $T=1404840 1473130 0 180 $X=1396100 $Y=1469190
X2231 13670 13652 12735 13626 13618 12811 24 13222 25 MXI4X1 $T=1404840 1546930 1 180 $X=1396100 $Y=1546678
X2232 13522 13614 12820 13625 13656 347 24 13250 25 MXI4X1 $T=1396560 1443610 1 0 $X=1396558 $Y=1439670
X2233 13716 13701 12820 13688 13671 386 24 13121 25 MXI4X1 $T=1409440 1421470 0 180 $X=1400700 $Y=1417530
X2234 13664 13623 12733 13609 13602 356 24 13252 25 MXI4X1 $T=1402540 1517410 1 0 $X=1402538 $Y=1513470
X2235 13716 13701 12729 13688 13671 12802 24 13227 25 MXI4X1 $T=1411740 1421470 1 180 $X=1403000 $Y=1421218
X2236 13665 13627 12729 13617 13604 367 24 13249 25 MXI4X1 $T=1404840 1369810 0 0 $X=1404838 $Y=1369558
X2237 13785 13761 12788 13749 13725 398 24 13144 25 MXI4X1 $T=1416340 1502650 0 180 $X=1407600 $Y=1498710
X2238 13775 13771 12790 13767 13753 365 24 13407 25 MXI4X1 $T=1418640 1399330 1 180 $X=1409900 $Y=1399078
X2239 13775 13771 12724 13767 13753 342 24 13223 25 MXI4X1 $T=1418640 1406710 1 180 $X=1409900 $Y=1406458
X2240 13791 13774 351 13768 13754 342 24 13358 25 MXI4X1 $T=1418640 1458370 0 180 $X=1409900 $Y=1454430
X2241 13785 13761 12718 13749 13725 364 24 13153 25 MXI4X1 $T=1418640 1495270 1 180 $X=1409900 $Y=1495018
X2242 460 459 354 465 467 367 24 13263 25 MXI4X1 $T=1410820 1355050 1 0 $X=1410818 $Y=1351110
X2243 13798 13780 12733 13770 13762 356 24 13128 25 MXI4X1 $T=1421400 1532170 1 180 $X=1412660 $Y=1531918
X2244 13702 13758 359 13779 13787 343 24 13242 25 MXI4X1 $T=1413580 1384570 0 0 $X=1413578 $Y=1384318
X2245 13791 13774 345 13768 13754 12828 24 13228 25 MXI4X1 $T=1422320 1450990 1 180 $X=1413580 $Y=1450738
X2246 13831 13756 12734 13786 13778 353 24 13232 25 MXI4X1 $T=1422320 1539550 1 180 $X=1413580 $Y=1539298
X2247 13702 13758 352 13779 13787 347 24 13377 25 MXI4X1 $T=1414040 1391950 1 0 $X=1414038 $Y=1388010
X2248 13831 13756 12735 13786 13778 12811 24 13115 25 MXI4X1 $T=1431060 1539550 1 180 $X=1422320 $Y=1539298
X2249 13865 13853 12788 13896 13925 383 24 13937 25 MXI4X1 $T=1426920 1473130 1 0 $X=1426918 $Y=1469190
X2250 13748 13823 12790 13895 13927 12828 24 13023 25 MXI4X1 $T=1427380 1421470 0 0 $X=1427378 $Y=1421218
X2251 13865 13853 12718 13896 13925 485 24 13941 25 MXI4X1 $T=1427380 1473130 0 0 $X=1427378 $Y=1472878
X2252 13871 13861 12735 13899 13854 398 24 13939 25 MXI4X1 $T=1427380 1510030 1 0 $X=1427378 $Y=1506090
X2253 13871 13861 12734 13899 13854 399 24 13892 25 MXI4X1 $T=1427380 1517410 1 0 $X=1427378 $Y=1513470
X2254 13748 13823 12724 13895 13927 342 24 13141 25 MXI4X1 $T=1430600 1428850 1 0 $X=1430598 $Y=1424910
X2255 13940 13954 12788 13964 13993 383 24 14050 25 MXI4X1 $T=1435660 1473130 1 0 $X=1435658 $Y=1469190
X2256 13971 13929 12734 13985 13970 353 24 13886 25 MXI4X1 $T=1444400 1495270 1 180 $X=1435660 $Y=1495018
X2257 13940 13954 12718 13964 13993 485 24 14052 25 MXI4X1 $T=1436120 1473130 0 0 $X=1436118 $Y=1472878
X2258 13949 13969 12788 13947 13958 382 24 14056 25 MXI4X1 $T=1437040 1443610 0 0 $X=1437038 $Y=1443358
X2259 13952 13965 444 13946 13953 492 24 14058 25 MXI4X1 $T=1437500 1384570 1 0 $X=1437498 $Y=1380630
X2260 13952 13965 442 13946 13953 374 24 14060 25 MXI4X1 $T=1437500 1384570 0 0 $X=1437498 $Y=1384318
X2261 13949 13969 12718 13947 13958 12802 24 14059 25 MXI4X1 $T=1437500 1443610 1 0 $X=1437498 $Y=1439670
X2262 13962 13982 12820 13976 13983 344 24 14063 25 MXI4X1 $T=1438420 1414090 0 0 $X=1438418 $Y=1413838
X2263 13971 13929 12735 13985 13970 12811 24 14114 25 MXI4X1 $T=1438880 1502650 1 0 $X=1438878 $Y=1498710
X2264 13962 13982 12729 13976 13983 485 24 14066 25 MXI4X1 $T=1439340 1414090 1 0 $X=1439338 $Y=1410150
X2265 14113 13950 12820 13989 13852 358 24 13998 25 MXI4X1 $T=1449920 1362430 1 180 $X=1441180 $Y=1362178
X2266 14031 14038 12734 14070 14115 343 24 14135 25 MXI4X1 $T=1444400 1517410 1 0 $X=1444398 $Y=1513470
X2267 14031 14038 12735 14070 14115 12811 24 14142 25 MXI4X1 $T=1444400 1524790 1 0 $X=1444398 $Y=1520850
X2268 14053 14062 12735 14071 14005 12811 24 14150 25 MXI4X1 $T=1444400 1546930 0 0 $X=1444398 $Y=1546678
X2269 14053 14062 12734 14071 14005 364 24 14182 25 MXI4X1 $T=1445780 1539550 0 0 $X=1445778 $Y=1539298
X2270 14262 14149 12820 14163 14159 401 24 14134 25 MXI4X1 $T=1460960 1436230 0 180 $X=1452220 $Y=1432290
X2271 14242 14227 12788 14160 14173 391 24 14139 25 MXI4X1 $T=1462340 1473130 1 180 $X=1453600 $Y=1472878
X2272 14113 13950 12729 13989 13852 485 24 14247 25 MXI4X1 $T=1454520 1369810 1 0 $X=1454518 $Y=1365870
X2273 14248 14184 12788 14192 14152 344 24 14122 25 MXI4X1 $T=1463260 1450990 0 180 $X=1454520 $Y=1447050
X2274 14251 14178 12735 14193 14177 12811 24 14153 25 MXI4X1 $T=1463260 1524790 0 180 $X=1454520 $Y=1520850
X2275 14145 14239 444 14195 14179 492 24 14124 25 MXI4X1 $T=1463720 1384570 0 180 $X=1454980 $Y=1380630
X2276 14242 14227 12718 14160 14173 485 24 14141 25 MXI4X1 $T=1464180 1480510 0 180 $X=1455440 $Y=1476570
X2277 14262 14149 12729 14163 14159 485 24 14162 25 MXI4X1 $T=1464640 1428850 0 180 $X=1455900 $Y=1424910
X2278 14248 14184 12718 14192 14152 485 24 14126 25 MXI4X1 $T=1465100 1443610 1 180 $X=1456360 $Y=1443358
X2279 14254 14246 12734 14175 14196 364 24 13978 25 MXI4X1 $T=1465100 1495270 1 180 $X=1456360 $Y=1495018
X2280 14314 14258 12820 14226 14232 391 24 14161 25 MXI4X1 $T=1466020 1414090 1 180 $X=1457280 $Y=1413838
X2281 14180 14237 12733 14250 14264 12811 24 14280 25 MXI4X1 $T=1459120 1539550 1 0 $X=1459118 $Y=1535610
X2282 14281 14266 12820 14257 14244 398 24 503 25 MXI4X1 $T=1467860 1362430 1 180 $X=1459120 $Y=1362178
X2283 14145 14239 442 14195 14179 386 24 14125 25 MXI4X1 $T=1459580 1384570 0 0 $X=1459578 $Y=1384318
X2284 14314 14258 12729 14226 14232 485 24 14224 25 MXI4X1 $T=1470620 1421470 0 180 $X=1461880 $Y=1417530
X2285 14180 14237 12810 14250 14264 384 24 14324 25 MXI4X1 $T=1462800 1532170 0 0 $X=1462798 $Y=1531918
X2286 14254 14246 12735 14175 14196 12811 24 14270 25 MXI4X1 $T=1463260 1502650 0 0 $X=1463258 $Y=1502398
X2287 14251 14178 12734 14193 14177 353 24 14240 25 MXI4X1 $T=1463260 1524790 1 0 $X=1463258 $Y=1520850
X2288 14281 14266 12729 14257 14244 492 24 14253 25 MXI4X1 $T=1472000 1369810 0 180 $X=1463260 $Y=1365870
X2289 14325 14272 12788 14276 14269 391 24 14147 25 MXI4X1 $T=1472000 1450990 0 180 $X=1463260 $Y=1447050
X2290 14327 14316 444 14279 14271 342 24 14151 25 MXI4X1 $T=1472460 1384570 0 180 $X=1463720 $Y=1380630
X2291 14325 14272 12718 14276 14269 485 24 14155 25 MXI4X1 $T=1473840 1443610 1 180 $X=1465100 $Y=1443358
X2292 14327 14316 442 14279 14271 382 24 14187 25 MXI4X1 $T=1474300 1391950 0 180 $X=1465560 $Y=1388010
X2293 511 514 352 14326 14338 358 24 14363 25 MXI4X1 $T=1468320 1362430 1 0 $X=1468318 $Y=1358490
X2294 511 514 359 14326 14338 343 24 14366 25 MXI4X1 $T=1469700 1362430 0 0 $X=1469698 $Y=1362178
X2295 14417 14381 13143 14324 14357 400 24 13302 25 MXI4X1 $T=1482120 1487890 0 180 $X=1473380 $Y=1483950
X2296 14378 14411 12733 14423 14432 12811 24 14433 25 MXI4X1 $T=1478900 1495270 0 0 $X=1478898 $Y=1495018
X2297 14414 14413 12790 14416 14448 12828 24 14462 25 MXI4X1 $T=1481200 1406710 0 0 $X=1481198 $Y=1406458
X2298 14378 14411 12810 14423 14432 525 24 14381 25 MXI4X1 $T=1481200 1487890 0 0 $X=1481198 $Y=1487638
X2299 14414 14413 12724 14416 14448 526 24 14464 25 MXI4X1 $T=1481660 1406710 1 0 $X=1481658 $Y=1402770
X2300 14335 14456 12724 14137 14512 342 24 14538 25 MXI4X1 $T=1486260 1384570 0 0 $X=1486258 $Y=1384318
X2301 14557 14534 12733 14520 14471 12811 24 14454 25 MXI4X1 $T=1496380 1502650 0 180 $X=1487640 $Y=1498710
X2302 14452 14458 345 14517 14529 12828 24 14565 25 MXI4X1 $T=1488560 1436230 1 0 $X=1488558 $Y=1432290
X2303 14452 14458 351 14517 14529 526 24 14569 25 MXI4X1 $T=1489020 1436230 0 0 $X=1489018 $Y=1435978
X2304 14461 14337 351 14465 14445 384 24 14562 25 MXI4X1 $T=1489020 1465750 0 0 $X=1489018 $Y=1465498
X2305 14453 14440 12733 14415 14420 356 24 14561 25 MXI4X1 $T=1489020 1517410 1 0 $X=1489018 $Y=1513470
X2306 14461 14337 345 14465 14445 356 24 14630 25 MXI4X1 $T=1489940 1465750 1 0 $X=1489938 $Y=1461810
X2307 14539 14558 12790 14540 14523 12828 24 14466 25 MXI4X1 $T=1498680 1406710 1 180 $X=1489940 $Y=1406458
X2308 14335 14456 12790 14137 14512 12828 24 14584 25 MXI4X1 $T=1490400 1391950 1 0 $X=1490398 $Y=1388010
X2309 14648 14363 30 13998 14527 396 24 13320 25 MXI4X1 $T=1499140 1362430 1 180 $X=1490400 $Y=1362178
X2310 14576 14466 107 14462 14528 396 24 13321 25 MXI4X1 $T=1499140 1406710 0 180 $X=1490400 $Y=1402770
X2311 14653 14563 345 14546 14530 356 24 14469 25 MXI4X1 $T=1499140 1495270 0 180 $X=1490400 $Y=1491330
X2312 14557 14534 12810 14520 14471 343 24 14357 25 MXI4X1 $T=1499140 1502650 1 180 $X=1490400 $Y=1502398
X2313 14522 14541 12733 14560 14571 356 24 14618 25 MXI4X1 $T=1492700 1517410 0 0 $X=1492698 $Y=1517158
X2314 14642 14590 12733 14460 14566 356 24 14533 25 MXI4X1 $T=1502820 1539550 0 180 $X=1494080 $Y=1535610
X2315 14635 536 334 14581 14575 533 24 14424 25 MXI4X1 $T=1504200 1369810 0 180 $X=1495460 $Y=1365870
X2316 14635 536 335 14581 14575 358 24 14527 25 MXI4X1 $T=1504660 1362430 0 180 $X=1495920 $Y=1358490
X2317 14568 14579 12790 14621 14631 12828 24 14637 25 MXI4X1 $T=1497760 1436230 1 0 $X=1497758 $Y=1432290
X2318 14568 14579 12724 14621 14631 526 24 14650 25 MXI4X1 $T=1497760 1436230 0 0 $X=1497758 $Y=1435978
X2319 14539 14558 12724 14540 14523 526 24 14636 25 MXI4X1 $T=1498680 1406710 0 0 $X=1498678 $Y=1406458
X2320 14655 14583 345 14628 14617 356 24 14587 25 MXI4X1 $T=1508800 1473130 0 180 $X=1500060 $Y=1469190
X2321 14743 14728 351 14683 14671 485 24 14627 25 MXI4X1 $T=1513400 1458370 1 180 $X=1504660 $Y=1458118
X2322 14644 14658 12724 14656 14697 526 24 14661 25 MXI4X1 $T=1505580 1384570 0 0 $X=1505578 $Y=1384318
X2323 14743 14728 345 14683 14671 356 24 14652 25 MXI4X1 $T=1515240 1458370 0 180 $X=1506500 $Y=1454430
X2324 14644 14658 12790 14656 14697 12828 24 14624 25 MXI4X1 $T=1509260 1391950 1 0 $X=1509258 $Y=1388010
X2325 14820 14775 541 14748 14753 12828 24 14646 25 MXI4X1 $T=1522140 1384570 0 180 $X=1513400 $Y=1380630
X2326 14823 14776 12790 14763 14754 12828 24 14528 25 MXI4X1 $T=1522140 1399330 1 180 $X=1513400 $Y=1399078
X2327 14669 14781 12790 14768 14757 12828 24 14663 25 MXI4X1 $T=1522600 1436230 0 180 $X=1513860 $Y=1432290
X2328 14820 14775 542 14748 14753 526 24 14696 25 MXI4X1 $T=1523060 1377190 1 180 $X=1514320 $Y=1376938
X2329 14823 14776 12724 14763 14754 526 24 14749 25 MXI4X1 $T=1523520 1406710 1 180 $X=1514780 $Y=1406458
X2330 14669 14781 12724 14768 14757 526 24 14752 25 MXI4X1 $T=1523980 1436230 1 180 $X=1515240 $Y=1435978
X2331 14786 14782 12733 14769 14759 356 24 14651 25 MXI4X1 $T=1520760 1517410 0 0 $X=1520758 $Y=1517158
X2332 14832 14777 345 14764 14755 356 24 14679 25 MXI4X1 $T=1540540 1495270 0 180 $X=1531800 $Y=1491330
X2333 80 24 32 25 CLKINVX12 $T=1116880 1369810 0 0 $X=1116878 $Y=1369558
X2334 10298 24 9741 25 CLKINVX12 $T=1138960 1480510 0 0 $X=1138958 $Y=1480258
X2335 10298 24 10663 25 CLKINVX12 $T=1211180 1465750 1 0 $X=1211178 $Y=1461810
X2336 10298 24 229 25 CLKINVX12 $T=1277420 1355050 0 0 $X=1277418 $Y=1354798
X2337 10298 24 12113 25 CLKINVX12 $T=1308700 1450990 0 0 $X=1308698 $Y=1450738
X2338 12720 24 11960 25 CLKINVX12 $T=1316060 1524790 0 0 $X=1316058 $Y=1524538
X2339 12720 24 13102 25 CLKINVX12 $T=1384600 1428850 0 0 $X=1384598 $Y=1428598
X2340 12720 24 13368 25 CLKINVX12 $T=1411280 1517410 1 0 $X=1411278 $Y=1513470
X2341 14144 24 466 25 CLKINVX12 $T=1452220 1377190 1 0 $X=1452218 $Y=1373250
X2342 14144 24 13766 25 CLKINVX12 $T=1453140 1473130 1 0 $X=1453138 $Y=1469190
X2343 14144 24 14256 25 CLKINVX12 $T=1508800 1510030 0 0 $X=1508798 $Y=1509778
X2344 14144 24 14370 25 CLKINVX12 $T=1523060 1428850 0 0 $X=1523058 $Y=1428598
X2345 13165 13159 12810 13145 13129 84 24 13278 25 MXI4XL $T=1359760 1532170 0 0 $X=1359758 $Y=1531918
X2346 13398 13375 12810 13322 13305 84 24 13237 25 MXI4XL $T=1375400 1517410 1 180 $X=1366660 $Y=1517158
X2347 13798 13780 12810 13770 13762 84 24 13253 25 MXI4XL $T=1419560 1532170 0 180 $X=1410820 $Y=1528230
X2348 14453 14440 12810 14415 14420 84 24 14376 25 MXI4XL $T=1487640 1517410 1 180 $X=1478900 $Y=1517158
X2349 14642 14590 12810 14460 14566 84 24 14547 25 MXI4XL $T=1505120 1532170 1 180 $X=1496380 $Y=1531918
X2350 14522 14541 12810 14560 14571 84 24 14535 25 MXI4XL $T=1497760 1524790 1 0 $X=1497758 $Y=1520850
X2351 14655 14583 351 14628 14617 84 24 14552 25 MXI4XL $T=1506500 1465750 1 180 $X=1497760 $Y=1465498
X2352 14653 14563 351 14546 14530 84 24 14545 25 MXI4XL $T=1507420 1487890 1 180 $X=1498680 $Y=1487638
X2353 14832 14777 351 14764 14755 84 24 14574 25 MXI4XL $T=1522140 1487890 1 180 $X=1513400 $Y=1487638
X2354 14786 14782 12810 14769 14759 84 24 14572 25 MXI4XL $T=1522600 1524790 0 180 $X=1513860 $Y=1520850
X2355 25 12489 309 12586 12581 24 12478 12602 12586 12113 296 12398 12581 12704 3961 ICV_29 $T=1299960 1428850 0 0 $X=1299958 $Y=1428598
X2356 25 12528 310 12587 12574 24 12478 12603 12587 12113 12404 12688 12574 12739 3961 ICV_29 $T=1299960 1436230 1 0 $X=1299958 $Y=1432290
X2357 25 12489 312 12589 12583 24 12597 12583 12610 12113 12404 12399 12599 12740 3961 ICV_29 $T=1299960 1465750 0 0 $X=1299958 $Y=1465498
X2358 25 12528 284 12568 12567 24 12370 12606 12568 11960 321 12342 12567 12698 3961 ICV_29 $T=1299960 1532170 1 0 $X=1299958 $Y=1528230
X2359 25 12726 310 12931 12917 24 289 12953 12962 229 380 12507 13056 13119 3961 ICV_29 $T=1334460 1391950 0 0 $X=1334458 $Y=1391698
X2360 25 12806 309 12933 12928 24 12478 12955 12933 12113 348 12688 12928 12966 3961 ICV_29 $T=1334460 1436230 0 0 $X=1334458 $Y=1435978
X2361 25 12726 274 12934 12929 24 12942 12949 12934 12113 381 12787 12929 13114 3961 ICV_29 $T=1334460 1450990 1 0 $X=1334458 $Y=1447050
X2362 25 12874 274 12935 12927 24 12597 12702 12935 12113 12641 12508 12927 13095 3961 ICV_29 $T=1334460 1450990 0 0 $X=1334458 $Y=1450738
X2363 25 12806 312 12919 12872 24 12597 12929 12919 12113 348 12560 12872 13106 3961 ICV_29 $T=1334460 1458370 1 0 $X=1334458 $Y=1454430
X2364 25 12874 284 12938 12873 24 12411 12956 12938 11960 12641 12974 12873 13026 3961 ICV_29 $T=1334460 1546930 0 0 $X=1334458 $Y=1546678
X2365 25 12806 274 12960 12955 24 12942 12907 12960 12113 348 12787 12955 13113 3961 ICV_29 $T=1336760 1443610 0 0 $X=1336758 $Y=1443358
X2366 25 413 13296 420 13360 24 366 13367 13389 13102 431 13476 13436 13489 3961 ICV_29 $T=1368960 1384570 1 0 $X=1368958 $Y=1380630
X2367 25 13517 312 13698 13696 24 13704 13712 13698 13102 454 12399 13696 13774 3961 ICV_29 $T=1403460 1465750 0 0 $X=1403458 $Y=1465498
X2368 25 489 471 14000 490 24 470 14041 14000 466 475 441 490 498 3961 ICV_29 $T=1437960 1355050 1 0 $X=1437958 $Y=1351110
X2369 25 488 471 14001 13994 24 470 13893 14001 466 480 441 13994 499 3961 ICV_29 $T=1437960 1355050 0 0 $X=1437958 $Y=1354798
X2370 25 13826 309 13975 14002 24 13659 14002 14045 466 495 12926 14138 14145 3961 ICV_29 $T=1437960 1399330 0 0 $X=1437958 $Y=1399078
X2371 25 14273 14356 14690 14692 24 14659 14689 14737 14370 524 13383 14760 14781 3961 ICV_29 $T=1506960 1421470 0 0 $X=1506958 $Y=1421218
X2372 12970 12932 30 13023 13038 43 25 24 13057 MX4X1 $T=1340900 1421470 0 0 $X=1340898 $Y=1421218
X2373 13063 12893 13107 13115 13135 393 25 24 13166 MX4X1 $T=1349640 1539550 0 0 $X=1349638 $Y=1539298
X2374 13054 12922 30 13121 13148 396 25 24 13181 MX4X1 $T=1350560 1421470 1 0 $X=1350558 $Y=1417530
X2375 13060 12813 13107 13128 13097 393 25 24 13177 MX4X1 $T=1351020 1532170 0 0 $X=1351018 $Y=1531918
X2376 13021 12817 30 13142 13163 43 25 24 13231 MX4X1 $T=1352400 1458370 0 0 $X=1352398 $Y=1458118
X2377 13100 12880 13107 13144 13164 393 25 24 13127 MX4X1 $T=1352400 1502650 1 0 $X=1352398 $Y=1498710
X2378 13116 12798 13143 13153 13172 400 25 24 13187 MX4X1 $T=1353320 1495270 0 0 $X=1353318 $Y=1495018
X2379 13111 12797 59 13219 13235 397 25 24 13245 MX4X1 $T=1358380 1465750 1 0 $X=1358378 $Y=1461810
X2380 13168 12891 13107 13220 13236 393 25 24 13229 MX4X1 $T=1358380 1487890 1 0 $X=1358378 $Y=1483950
X2381 13059 12845 13143 13221 13237 400 25 24 13122 MX4X1 $T=1358380 1510030 0 0 $X=1358378 $Y=1509778
X2382 13169 12899 13107 13222 13239 393 25 24 13247 MX4X1 $T=1358380 1539550 0 0 $X=1358378 $Y=1539298
X2383 13161 12807 59 13223 13243 397 25 24 13234 MX4X1 $T=1358840 1406710 1 0 $X=1358838 $Y=1402770
X2384 13171 12837 13143 13224 13246 400 25 24 13276 MX4X1 $T=1358840 1487890 0 0 $X=1358838 $Y=1487638
X2385 13130 12814 403 13227 13255 397 25 24 13226 MX4X1 $T=1359760 1421470 1 0 $X=1359758 $Y=1417530
X2386 13178 12890 30 13228 13256 410 25 24 13295 MX4X1 $T=1359760 1450990 0 0 $X=1359758 $Y=1450738
X2387 13098 12816 13143 13232 13262 400 25 24 13238 MX4X1 $T=1360220 1546930 1 0 $X=1360218 $Y=1542990
X2388 13189 12959 404 13242 13271 60 25 24 13296 MX4X1 $T=1361140 1384570 0 0 $X=1361138 $Y=1384318
X2389 13216 13033 405 13249 13274 412 25 24 13306 MX4X1 $T=1361600 1377190 1 0 $X=1361598 $Y=1373250
X2390 13217 12918 107 13250 13275 393 25 24 13288 MX4X1 $T=1361600 1443610 0 0 $X=1361598 $Y=1443358
X2391 13031 12923 13107 13252 13277 393 25 24 13304 MX4X1 $T=1361600 1517410 1 0 $X=1361598 $Y=1513470
X2392 13218 12892 13143 13253 13278 400 25 24 13230 MX4X1 $T=1361600 1532170 1 0 $X=1361598 $Y=1528230
X2393 13175 12915 405 13263 13293 412 25 24 419 MX4X1 $T=1362980 1355050 1 0 $X=1362978 $Y=1351110
X2394 13185 12903 59 13358 13393 397 25 24 13349 MX4X1 $T=1368960 1458370 1 0 $X=1368958 $Y=1454430
X2395 13273 12882 13143 13372 13392 412 25 24 13371 MX4X1 $T=1369880 1450990 1 0 $X=1369878 $Y=1447050
X2396 13268 12905 428 13377 13404 410 25 24 13390 MX4X1 $T=1370340 1391950 1 0 $X=1370338 $Y=1388010
X2397 13978 13892 13143 13886 13876 400 25 24 13248 MX4X1 $T=1432440 1495270 0 180 $X=1423700 $Y=1491330
X2398 14139 13937 13107 14050 14065 393 25 24 13285 MX4X1 $T=1453140 1473130 0 180 $X=1444400 $Y=1469190
X2399 14141 13941 13143 14052 14067 400 25 24 13386 MX4X1 $T=1453600 1473130 1 180 $X=1444860 $Y=1472878
X2400 14147 14056 433 14122 14072 43 25 24 13314 MX4X1 $T=1454520 1443610 1 180 $X=1445780 $Y=1443358
X2401 14151 14058 404 14124 14073 60 25 24 13360 MX4X1 $T=1454980 1384570 0 180 $X=1446240 $Y=1380630
X2402 14187 14060 428 14125 14074 410 25 24 13426 MX4X1 $T=1454980 1384570 1 180 $X=1446240 $Y=1384318
X2403 14155 14059 403 14126 14075 412 25 24 13400 MX4X1 $T=1454980 1443610 0 180 $X=1446240 $Y=1439670
X2404 14161 14063 30 14134 14117 410 25 24 13301 MX4X1 $T=1455900 1414090 1 180 $X=1447160 $Y=1413838
X2405 14153 14150 13107 14142 14127 393 25 24 13259 MX4X1 $T=1457280 1517410 1 180 $X=1448540 $Y=1517158
X2406 14224 14066 403 14162 14146 400 25 24 13257 MX4X1 $T=1460040 1414090 0 180 $X=1451300 $Y=1410150
X2407 14240 14182 13143 14135 14165 400 25 24 13265 MX4X1 $T=1461880 1517410 0 180 $X=1453140 $Y=1513470
X2408 14253 507 405 506 14183 412 25 24 500 MX4X1 $T=1464640 1355050 0 180 $X=1455900 $Y=1351110
X2409 14270 13939 13107 14114 14185 393 25 24 13157 MX4X1 $T=1464640 1510030 0 180 $X=1455900 $Y=1506090
X2410 14424 14247 405 14366 14354 412 25 24 13394 MX4X1 $T=1482120 1369810 0 180 $X=1473380 $Y=1365870
X2411 14454 14280 13107 14433 14418 393 25 24 13286 MX4X1 $T=1487640 1502650 0 180 $X=1478900 $Y=1498710
X2412 14572 14547 13143 14535 14516 400 25 24 13291 MX4X1 $T=1497760 1524790 0 180 $X=1489020 $Y=1520850
X2413 14574 14376 13143 14545 14521 400 25 24 13150 MX4X1 $T=1498680 1487890 1 180 $X=1489940 $Y=1487638
X2414 14627 14562 59 14552 14524 397 25 24 13281 MX4X1 $T=1499140 1458370 1 180 $X=1490400 $Y=1458118
X2415 14679 14561 13107 14469 14577 393 25 24 13374 MX4X1 $T=1505120 1495270 1 180 $X=1496380 $Y=1495018
X2416 14646 14584 433 14624 14582 43 25 24 13104 MX4X1 $T=1505580 1384570 1 180 $X=1496840 $Y=1384318
X2417 14652 14630 30 14587 14588 43 25 24 13284 MX4X1 $T=1506500 1458370 0 180 $X=1497760 $Y=1454430
X2418 14651 14533 13107 14618 14589 393 25 24 13251 MX4X1 $T=1506500 1517410 0 180 $X=1497760 $Y=1513470
X2419 14749 14464 59 14636 14625 397 25 24 13269 MX4X1 $T=1507880 1406710 0 180 $X=1499140 $Y=1402770
X2420 14663 14565 30 14637 14626 43 25 24 13363 MX4X1 $T=1507880 1428850 1 180 $X=1499140 $Y=1428598
X2421 14696 14538 59 14661 14643 397 25 24 13233 MX4X1 $T=1511100 1384570 0 180 $X=1502360 $Y=1380630
X2422 14752 14569 59 14650 14681 397 25 24 13403 MX4X1 $T=1515240 1436230 1 180 $X=1506500 $Y=1435978
X2423 44 13127 394 13157 24 25 MXI2X2 $T=1352860 1502650 0 0 $X=1352858 $Y=1502398
X2424 44 13166 11898 13259 24 25 MXI2X2 $T=1357920 1510030 1 0 $X=1357918 $Y=1506090
X2425 44 13229 406 13285 24 25 MXI2X2 $T=1361600 1473130 1 0 $X=1361598 $Y=1469190
X2426 417 13314 416 13288 24 25 MXI2X2 $T=1372640 1443610 0 180 $X=1368040 $Y=1439670
X2427 44 13304 421 13374 24 25 MXI2X2 $T=1368960 1495270 1 0 $X=1368958 $Y=1491330
X2428 414 13390 432 13426 24 25 MXI2X2 $T=1373100 1384570 0 0 $X=1373098 $Y=1384318
X2429 26 27 25 24 INVX12 $T=747960 1465750 1 0 $X=747958 $Y=1461810
X2430 7872 28 25 24 INVX12 $T=757160 1495270 1 0 $X=757158 $Y=1491330
X2431 10914 161 25 24 INVX12 $T=1190480 1384570 1 180 $X=1186800 $Y=1384318
X2432 11017 160 25 24 INVX12 $T=1192320 1406710 0 180 $X=1188640 $Y=1402770
X2433 11166 175 25 24 INVX12 $T=1213480 1436230 0 0 $X=1213478 $Y=1435978
X2434 11311 201 25 24 INVX12 $T=1223140 1443610 1 180 $X=1219460 $Y=1443358
X2435 11438 197 25 24 INVX12 $T=1228200 1473130 0 180 $X=1224520 $Y=1469190
X2436 11480 208 25 24 INVX12 $T=1231880 1487890 1 0 $X=1231878 $Y=1483950
X2437 11632 217 25 24 INVX12 $T=1244300 1487890 0 180 $X=1240620 $Y=1483950
X2438 11356 245 25 24 INVX12 $T=1252120 1517410 0 0 $X=1252118 $Y=1517158
X2439 11954 241 25 24 INVX12 $T=1259020 1436230 1 180 $X=1255340 $Y=1435978
X2440 12207 269 25 24 INVX12 $T=1277880 1510030 1 0 $X=1277878 $Y=1506090
X2441 12205 272 25 24 INVX12 $T=1284320 1436230 0 0 $X=1284318 $Y=1435978
X2442 11777 290 25 24 INVX12 $T=1284320 1473130 1 0 $X=1284318 $Y=1469190
X2443 12244 286 25 24 INVX12 $T=1284320 1495270 0 0 $X=1284318 $Y=1495018
X2444 11206 292 25 24 INVX12 $T=1284780 1421470 1 0 $X=1284778 $Y=1417530
X2445 11902 281 25 24 INVX12 $T=1286620 1458370 0 0 $X=1286618 $Y=1458118
X2446 12115 362 25 24 INVX12 $T=1327560 1487890 1 0 $X=1327558 $Y=1483950
X2447 12056 370 25 24 INVX12 $T=1334460 1480510 1 0 $X=1334458 $Y=1476570
X2448 12243 436 25 24 INVX12 $T=1371260 1480510 1 0 $X=1371258 $Y=1476570
X2449 10760 10733 10716 25 24 10713 CLKMX2X2 $T=1176680 1414090 1 180 $X=1173000 $Y=1413838
X2450 10760 10780 10721 25 24 10717 CLKMX2X2 $T=1177600 1421470 0 0 $X=1177598 $Y=1421218
X2451 10760 10946 10897 25 24 10807 CLKMX2X2 $T=1188640 1436230 1 180 $X=1184960 $Y=1435978
X2452 10760 10969 10794 25 24 10761 CLKMX2X2 $T=1194160 1428850 1 180 $X=1190480 $Y=1428598
X2453 10760 11108 11079 25 24 10944 CLKMX2X2 $T=1200140 1399330 1 180 $X=1196460 $Y=1399078
X2454 10760 11119 11075 25 24 10950 CLKMX2X2 $T=1200600 1450990 1 180 $X=1196920 $Y=1450738
X2455 10760 11199 11163 25 24 11029 CLKMX2X2 $T=1205660 1473130 0 180 $X=1201980 $Y=1469190
X2456 162 182 11175 25 24 11299 CLKMX2X2 $T=1207040 1362430 0 0 $X=1207038 $Y=1362178
X2457 10952 11358 11308 25 24 11167 CLKMX2X2 $T=1217620 1480510 0 180 $X=1213940 $Y=1476570
X2458 162 194 11324 25 24 11371 CLKMX2X2 $T=1214860 1362430 0 0 $X=1214858 $Y=1362178
X2459 10952 11338 11364 25 24 11076 CLKMX2X2 $T=1214860 1502650 0 0 $X=1214858 $Y=1502398
X2460 10952 11345 11369 25 24 11198 CLKMX2X2 $T=1215320 1524790 0 0 $X=1215318 $Y=1524538
X2461 10952 11382 11430 25 24 11195 CLKMX2X2 $T=1219000 1495270 0 0 $X=1218998 $Y=1495018
X2462 162 204 11394 25 24 11507 CLKMX2X2 $T=1224520 1362430 1 0 $X=1224518 $Y=1358490
X2463 10952 11510 11463 25 24 11476 CLKMX2X2 $T=1228660 1517410 0 180 $X=1224980 $Y=1513470
X2464 162 209 11594 25 24 11638 CLKMX2X2 $T=1230500 1377190 1 0 $X=1230498 $Y=1373250
X2465 10760 11607 11583 25 24 11449 CLKMX2X2 $T=1234640 1414090 1 180 $X=1230960 $Y=1413838
X2466 10952 11597 11620 25 24 11658 CLKMX2X2 $T=1232340 1517410 0 0 $X=1232338 $Y=1517158
X2467 162 212 11641 25 24 11645 CLKMX2X2 $T=1233720 1369810 1 0 $X=1233718 $Y=1365870
X2468 162 215 11586 25 24 11667 CLKMX2X2 $T=1235560 1355050 1 0 $X=1235558 $Y=1351110
X2469 10760 11698 11736 25 24 11668 CLKMX2X2 $T=1241540 1406710 0 0 $X=1241538 $Y=1406458
X2470 10952 11742 11744 25 24 11532 CLKMX2X2 $T=1245680 1517410 1 180 $X=1242000 $Y=1517158
X2471 162 228 11807 25 24 11875 CLKMX2X2 $T=1246600 1362430 0 0 $X=1246598 $Y=1362178
X2472 157 232 11898 25 24 238 CLKMX2X2 $T=1249360 1355050 1 0 $X=1249358 $Y=1351110
X2473 10760 11876 235 25 24 11905 CLKMX2X2 $T=1249360 1406710 1 0 $X=1249358 $Y=1402770
X2474 157 237 11882 25 24 11773 CLKMX2X2 $T=1253040 1377190 1 180 $X=1249360 $Y=1376938
X2475 157 242 11947 25 24 225 CLKMX2X2 $T=1254880 1384570 0 0 $X=1254878 $Y=1384318
X2476 10952 11966 11948 25 24 11893 CLKMX2X2 $T=1260400 1517410 1 180 $X=1256720 $Y=1517158
X2477 157 247 12018 25 24 251 CLKMX2X2 $T=1258100 1355050 1 0 $X=1258098 $Y=1351110
X2478 157 226 12020 25 24 11899 CLKMX2X2 $T=1258560 1384570 1 0 $X=1258558 $Y=1380630
X2479 157 239 12021 25 24 253 CLKMX2X2 $T=1258560 1391950 1 0 $X=1258558 $Y=1388010
X2480 11123 12016 12035 25 24 11873 CLKMX2X2 $T=1259940 1421470 0 0 $X=1259938 $Y=1421218
X2481 157 244 12081 25 24 11798 CLKMX2X2 $T=1264540 1391950 1 0 $X=1264538 $Y=1388010
X2482 157 246 12084 25 24 257 CLKMX2X2 $T=1265000 1384570 1 0 $X=1264998 $Y=1380630
X2483 157 254 12093 25 24 11924 CLKMX2X2 $T=1265460 1384570 0 0 $X=1265458 $Y=1384318
X2484 10952 12092 12075 25 24 11943 CLKMX2X2 $T=1269140 1524790 0 180 $X=1265460 $Y=1520850
X2485 102 243 12193 25 24 223 CLKMX2X2 $T=1270980 1384570 1 0 $X=1270978 $Y=1380630
X2486 10952 12200 12222 25 24 12103 CLKMX2X2 $T=1273740 1524790 0 0 $X=1273738 $Y=1524538
X2487 102 259 12237 25 24 11877 CLKMX2X2 $T=1276040 1377190 1 0 $X=1276038 $Y=1373250
X2488 10952 12247 12201 25 24 12099 CLKMX2X2 $T=1280180 1524790 0 180 $X=1276500 $Y=1520850
X2489 157 252 12245 25 24 249 CLKMX2X2 $T=1276960 1384570 1 0 $X=1276958 $Y=1380630
X2490 157 255 12251 25 24 267 CLKMX2X2 $T=1277420 1355050 1 0 $X=1277418 $Y=1351110
X2491 102 261 12252 25 24 11894 CLKMX2X2 $T=1277420 1428850 0 0 $X=1277418 $Y=1428598
X2492 102 273 12351 25 24 11675 CLKMX2X2 $T=1282020 1428850 0 0 $X=1282018 $Y=1428598
X2493 73 12518 10507 25 24 12580 CLKMX2X2 $T=1299040 1362430 1 0 $X=1299038 $Y=1358490
X2494 414 13184 13320 25 24 424 CLKMX2X2 $T=1368960 1362430 0 0 $X=1368958 $Y=1362178
X2495 44 13297 13321 25 24 425 CLKMX2X2 $T=1368960 1406710 1 0 $X=1368958 $Y=1402770
X2496 413 13352 13302 25 24 12093 CLKMX2X2 $T=1372640 1480510 1 180 $X=1368960 $Y=1480258
X2497 10005 24 25 10382 INVX2 $T=1145860 1369810 1 0 $X=1145858 $Y=1365870
X2498 10126 24 25 9920 INVX2 $T=1146320 1399330 0 0 $X=1146318 $Y=1399078
X2499 10735 24 25 10628 INVX2 $T=1173920 1377190 1 0 $X=1173918 $Y=1373250
X2500 11383 24 25 409 INVX2 $T=1362060 1377190 0 0 $X=1362058 $Y=1376938
X2501 11794 24 187 25 CLKINVX8 $T=1359760 1355050 1 0 $X=1359758 $Y=1351110
X2502 13058 12971 59 13141 13162 397 25 24 13188 MX4XL $T=1352400 1428850 1 0 $X=1352398 $Y=1424910
X2503 10614 25 10583 10502 24 NOR2XL $T=1164260 1473130 1 180 $X=1162880 $Y=1472878
X2504 134 25 131 10644 24 NOR2XL $T=1165640 1362430 0 0 $X=1165638 $Y=1362178
X2505 10623 25 131 10736 24 NOR2XL $T=1170240 1362430 0 0 $X=1170238 $Y=1362178
X2506 10676 25 10628 10756 24 NOR2XL $T=1173920 1473130 1 0 $X=1173918 $Y=1469190
X2507 10599 25 10773 10729 24 NOR2XL $T=1176680 1517410 1 180 $X=1175300 $Y=1517158
X2508 10811 25 10599 10851 24 NOR2XL $T=1179440 1524790 0 0 $X=1179438 $Y=1524538
X2509 10672 25 10628 10864 24 NOR2XL $T=1179900 1473130 1 0 $X=1179898 $Y=1469190
X2510 10599 25 10866 10769 24 NOR2XL $T=1182200 1502650 1 180 $X=1180820 $Y=1502398
X2511 10599 25 10867 10633 24 NOR2XL $T=1182200 1517410 0 180 $X=1180820 $Y=1513470
X2512 10599 25 10868 10771 24 NOR2XL $T=1182200 1517410 1 180 $X=1180820 $Y=1517158
X2513 10947 25 10867 11070 24 NOR2XL $T=1192320 1510030 0 0 $X=1192318 $Y=1509778
X2514 12201 25 10743 12170 24 NOR2XL $T=1272360 1458370 1 180 $X=1270980 $Y=1458118
X2515 77 25 68 12901 24 NOR2XL $T=1330780 1362430 1 0 $X=1330778 $Y=1358490
X2516 77 25 12812 12916 24 NOR2XL $T=1331700 1362430 0 0 $X=1331698 $Y=1362178
X2517 10947 10599 25 24 10770 NOR2BXL $T=1182660 1510030 0 180 $X=1180820 $Y=1506090
X2518 77 12812 25 24 12736 NOR2BXL $T=1326180 1362430 1 180 $X=1324340 $Y=1362178
X2519 77 68 25 24 12884 NOR2BXL $T=1331240 1369810 1 0 $X=1331238 $Y=1365870
X2520 10126 92 24 25 INVX3 $T=1139420 1414090 1 0 $X=1139418 $Y=1410150
X2521 104 82 24 25 INVX3 $T=1140800 1377190 1 0 $X=1140798 $Y=1373250
X2522 10333 107 24 25 INVX3 $T=1144940 1384570 1 0 $X=1144938 $Y=1380630
X2523 39 10245 24 25 INVX3 $T=1294440 1443610 1 0 $X=1294438 $Y=1439670
X2524 10382 127 24 25 INVX3 $T=1323420 1369810 0 0 $X=1323418 $Y=1369558
X2525 328 24 12720 25 CLKBUFX16 $T=1311460 1414090 1 0 $X=1311458 $Y=1410150
X2526 328 24 80 25 CLKBUFX16 $T=1315140 1406710 0 0 $X=1315138 $Y=1406458
X2527 10371 24 10274 10251 25 NAND2XL $T=1146320 1480510 0 180 $X=1144940 $Y=1476570
X2528 10389 24 10460 10465 25 NAND2XL $T=1150000 1487890 1 0 $X=1149998 $Y=1483950
X2529 148 24 10806 10875 25 NAND2XL $T=1178520 1369810 0 0 $X=1178518 $Y=1369558
X2530 10963 24 156 11078 25 NAND2XL $T=1191400 1369810 1 0 $X=1191398 $Y=1365870
X2531 10935 24 10953 10963 25 NAND2XL $T=1192780 1362430 0 180 $X=1191400 $Y=1358490
X2532 10970 24 10817 10951 25 NAND2XL $T=1194160 1487890 0 180 $X=1192780 $Y=1483950
X2533 11328 24 11357 11391 25 NAND2XL $T=1216700 1369810 1 0 $X=1216698 $Y=1365870
X2534 206 24 207 11525 25 NAND2XL $T=1226820 1355050 1 0 $X=1226818 $Y=1351110
X2535 11486 24 10778 11522 25 NAND2XL $T=1226820 1384570 1 0 $X=1226818 $Y=1380630
X2536 11364 24 11051 11534 25 NAND2XL $T=1229580 1443610 0 0 $X=1229578 $Y=1443358
X2537 11463 24 11063 11593 25 NAND2XL $T=1231420 1473130 0 0 $X=1231418 $Y=1472878
X2538 220 24 219 11652 25 NAND2XL $T=1242000 1355050 0 180 $X=1240620 $Y=1351110
X2539 11649 24 11735 11684 25 NAND2XL $T=1244300 1436230 0 180 $X=1242920 $Y=1432290
X2540 10137 24 10033 12671 25 NAND2XL $T=1311920 1369810 1 0 $X=1311918 $Y=1365870
X2541 12330 274 24 12114 12347 25 12357 12377 OAI221XL $T=1282480 1450990 1 0 $X=1282478 $Y=1447050
X2542 279 280 24 12355 12364 25 12368 12378 OAI221XL $T=1283860 1369810 1 0 $X=1283858 $Y=1365870
X2543 12330 284 24 12318 12347 25 12387 12389 OAI221XL $T=1285240 1517410 0 0 $X=1285238 $Y=1517158
X2544 279 295 24 12412 12364 25 12405 12397 OAI221XL $T=1292140 1384570 1 180 $X=1288920 $Y=1384318
X2545 12330 308 24 12472 12347 25 12473 12468 OAI221XL $T=1295820 1517410 0 180 $X=1292600 $Y=1513470
X2546 12330 299 24 12481 12347 25 12358 12501 OAI221XL $T=1293520 1428850 1 0 $X=1293518 $Y=1424910
X2547 12330 300 24 12465 12347 25 12471 12502 OAI221XL $T=1293520 1465750 0 0 $X=1293518 $Y=1465498
X2548 12330 298 24 12386 12347 25 12487 12523 OAI221XL $T=1293520 1495270 0 0 $X=1293518 $Y=1495018
X2549 12330 312 24 12317 12347 25 12480 12464 OAI221XL $T=1297200 1473130 0 180 $X=1293980 $Y=1469190
X2550 12330 305 24 12466 12347 25 12512 12503 OAI221XL $T=1295360 1487890 1 0 $X=1295358 $Y=1483950
X2551 12330 310 24 12356 12347 25 12566 12527 OAI221XL $T=1299500 1414090 0 0 $X=1299498 $Y=1413838
X2552 279 311 24 12509 12347 25 12570 12585 OAI221XL $T=1299960 1384570 1 0 $X=1299958 $Y=1380630
X2553 12330 309 24 12510 12347 25 12572 12588 OAI221XL $T=1299960 1436230 0 0 $X=1299958 $Y=1435978
X2554 12330 313 24 12504 12347 25 12524 12592 OAI221XL $T=1299960 1502650 1 0 $X=1299958 $Y=1498710
X2555 12330 301 24 12519 12347 25 12613 12632 OAI221XL $T=1303640 1517410 1 0 $X=1303638 $Y=1513470
X2556 101 12189 24 12671 12673 25 12253 12636 OAI221XL $T=1310080 1384570 0 0 $X=1310078 $Y=1384318
X2557 12329 275 12336 277 24 25 12368 OA22X1 $T=1282480 1362430 0 0 $X=1282478 $Y=1362178
X2558 12349 275 12365 277 24 25 12405 OA22X1 $T=1284780 1391950 1 0 $X=1284778 $Y=1388010
X2559 12353 12253 11922 12366 24 25 12471 OA22X1 $T=1284780 1465750 0 0 $X=1284778 $Y=1465498
X2560 12384 12253 12369 12366 24 25 12358 OA22X1 $T=1287540 1428850 0 180 $X=1284780 $Y=1424910
X2561 12206 12253 11470 12366 24 25 12473 OA22X1 $T=1288460 1524790 1 0 $X=1288458 $Y=1520850
X2562 12467 12253 12479 12366 24 25 12357 OA22X1 $T=1295820 1450990 1 180 $X=1293060 $Y=1450738
X2563 12415 12253 12486 12366 24 25 12512 OA22X1 $T=1294900 1487890 0 0 $X=1294898 $Y=1487638
X2564 12416 12253 12488 12366 24 25 12524 OA22X1 $T=1294900 1502650 1 0 $X=1294898 $Y=1498710
X2565 12505 12253 12474 12366 24 25 12387 OA22X1 $T=1297660 1524790 0 180 $X=1294900 $Y=1520850
X2566 12490 12253 12413 12366 24 25 12566 OA22X1 $T=1299960 1421470 1 0 $X=1299958 $Y=1417530
X2567 12584 12253 12564 12366 24 25 12487 OA22X1 $T=1302720 1495270 1 180 $X=1299960 $Y=1495018
X2568 12482 12253 12496 12366 24 25 12480 OA22X1 $T=1301340 1473130 1 0 $X=1301338 $Y=1469190
X2569 12565 12253 12382 12366 24 25 12613 OA22X1 $T=1302260 1517410 0 0 $X=1302258 $Y=1517158
X2570 12511 12253 12573 12366 24 25 12572 OA22X1 $T=1303640 1443610 1 0 $X=1303638 $Y=1439670
X2571 12608 12253 12166 277 24 25 12570 OA22X1 $T=1306400 1391950 1 0 $X=1306398 $Y=1388010
X2572 12614 275 323 277 24 25 326 OA22X1 $T=1307320 1355050 1 0 $X=1307318 $Y=1351110
X2573 9830 9682 36 24 9805 25 9753 AO22X1 $T=1095260 1436230 0 180 $X=1092500 $Y=1432290
X2574 9830 9674 40 24 9805 25 9747 AO22X1 $T=1097100 1428850 1 180 $X=1094340 $Y=1428598
X2575 9830 9678 42 24 9805 25 9749 AO22X1 $T=1097560 1450990 0 180 $X=1094800 $Y=1447050
X2576 9830 9902 48 24 9805 25 9755 AO22X1 $T=1100320 1450990 1 180 $X=1097560 $Y=1450738
X2577 9830 9823 52 24 9805 25 9923 AO22X1 $T=1103080 1428850 0 0 $X=1103078 $Y=1428598
X2578 9830 9934 56 24 9805 25 9921 AO22X1 $T=1106760 1480510 0 180 $X=1104000 $Y=1476570
X2579 9830 9994 63 24 9805 25 9806 AO22X1 $T=1111820 1443610 1 180 $X=1109060 $Y=1443358
X2580 9830 9993 64 24 9805 25 10027 AO22X1 $T=1109520 1480510 0 0 $X=1109518 $Y=1480258
X2581 9830 10004 67 24 9805 25 9835 AO22X1 $T=1112740 1465750 0 180 $X=1109980 $Y=1461810
X2582 9830 10013 69 24 9805 25 9991 AO22X1 $T=1114580 1458370 1 180 $X=1111820 $Y=1458118
X2583 9830 10034 71 24 9805 25 10057 AO22X1 $T=1113660 1487890 0 0 $X=1113658 $Y=1487638
X2584 9830 10067 78 24 9805 25 10010 AO22X1 $T=1118720 1465750 0 180 $X=1115960 $Y=1461810
X2585 10146 10124 82 24 58 25 10058 AO22X1 $T=1122860 1428850 1 180 $X=1120100 $Y=1428598
X2586 10146 10143 82 24 9745 25 9951 AO22X1 $T=1124700 1436230 0 180 $X=1121940 $Y=1432290
X2587 9830 10006 87 24 9805 25 10128 AO22X1 $T=1125160 1473130 1 180 $X=1122400 $Y=1472878
X2588 9830 10180 95 24 9805 25 10118 AO22X1 $T=1131600 1495270 1 180 $X=1128840 $Y=1495018
X2589 10146 10255 82 24 97 25 10229 AO22X1 $T=1136660 1428850 1 180 $X=1133900 $Y=1428598
X2590 10146 10270 82 24 10246 25 10357 AO22X1 $T=1142640 1414090 1 0 $X=1142638 $Y=1410150
X2591 10146 10270 82 24 10367 25 10394 AO22X1 $T=1144020 1428850 1 0 $X=1144018 $Y=1424910
X2592 10387 10369 108 24 9805 25 10175 AO22X1 $T=1146780 1517410 0 180 $X=1144020 $Y=1513470
X2593 10146 10375 82 24 10355 25 10235 AO22X1 $T=1147700 1421470 1 180 $X=1144940 $Y=1421218
X2594 9830 10474 117 24 9805 25 10368 AO22X1 $T=1153220 1502650 0 180 $X=1150460 $Y=1498710
X2595 10387 10488 122 24 10578 25 10476 AO22X1 $T=1162420 1502650 0 180 $X=1159660 $Y=1498710
X2596 9830 10636 132 24 10578 25 10611 AO22X1 $T=1166560 1487890 0 180 $X=1163800 $Y=1483950
X2597 10387 10568 143 24 10578 25 10448 AO22X1 $T=1171620 1510030 0 0 $X=1171618 $Y=1509778
X2598 165 10615 10964 24 10505 25 10947 AO22X1 $T=1191860 1510030 0 180 $X=1189100 $Y=1506090
X2599 162 163 10883 24 164 25 11034 AO22X1 $T=1189560 1355050 1 0 $X=1189558 $Y=1351110
X2600 162 169 10759 24 10279 25 11074 AO22X1 $T=1194620 1362430 0 0 $X=1194618 $Y=1362178
X2601 162 172 11096 24 164 25 11124 AO22X1 $T=1197840 1369810 0 0 $X=1197838 $Y=1369558
X2602 162 185 10927 24 164 25 11182 AO22X1 $T=1209340 1369810 1 180 $X=1206580 $Y=1369558
X2603 162 188 11116 24 164 25 11221 AO22X1 $T=1210260 1377190 1 180 $X=1207500 $Y=1376938
X2604 162 205 11432 24 10279 25 11453 AO22X1 $T=1226820 1362430 1 180 $X=1224060 $Y=1362178
X2605 162 213 11490 24 164 25 11545 AO22X1 $T=1235560 1384570 0 180 $X=1232800 $Y=1380630
X2606 162 216 11578 24 164 25 11584 AO22X1 $T=1236940 1384570 1 180 $X=1234180 $Y=1384318
X2607 11179 11675 11669 24 10279 25 11655 AO22X1 $T=1240620 1458370 0 180 $X=1237860 $Y=1454430
X2608 162 222 11749 24 164 25 11625 AO22X1 $T=1244760 1399330 1 180 $X=1242000 $Y=1399078
X2609 11179 223 11677 24 164 25 11654 AO22X1 $T=1244760 1450990 0 180 $X=1242000 $Y=1447050
X2610 11179 11798 11802 24 164 25 11889 AO22X1 $T=1247060 1450990 1 0 $X=1247058 $Y=1447050
X2611 11179 11877 11699 24 164 25 11589 AO22X1 $T=1250740 1428850 1 180 $X=1247980 $Y=1428598
X2612 11179 11773 11869 24 164 25 11921 AO22X1 $T=1248440 1428850 1 0 $X=1248438 $Y=1424910
X2613 11179 11894 11890 24 10279 25 11612 AO22X1 $T=1252120 1458370 0 180 $X=1249360 $Y=1454430
X2614 11179 249 11967 24 164 25 11883 AO22X1 $T=1260860 1450990 1 180 $X=1258100 $Y=1450738
X2615 11179 11899 12061 24 164 25 12068 AO22X1 $T=1264080 1458370 1 0 $X=1264078 $Y=1454430
X2616 11179 11924 12070 24 10279 25 12022 AO22X1 $T=1267760 1473130 0 180 $X=1265000 $Y=1469190
X2617 11179 225 12071 24 164 25 12172 AO22X1 $T=1265460 1436230 1 0 $X=1265458 $Y=1432290
X2618 11179 253 12072 24 164 25 12169 AO22X1 $T=1265460 1458370 0 0 $X=1265458 $Y=1458118
X2619 11179 257 12086 24 10279 25 12069 AO22X1 $T=1268680 1465750 1 180 $X=1265920 $Y=1465498
X2620 276 11662 283 24 12348 25 12407 AO22X1 $T=1283400 1377190 0 0 $X=1283398 $Y=1376938
X2621 276 11744 283 24 12177 25 12393 AO22X1 $T=1283400 1487890 0 0 $X=1283398 $Y=1487638
X2622 276 12075 283 24 12361 25 12340 AO22X1 $T=1283400 1502650 1 0 $X=1283398 $Y=1498710
X2623 276 12187 285 24 12102 25 12236 AO22X1 $T=1286160 1443610 1 180 $X=1283400 $Y=1443358
X2624 276 12201 283 24 12339 25 12337 AO22X1 $T=1286160 1473130 1 180 $X=1283400 $Y=1472878
X2625 276 11463 285 24 12232 25 12406 AO22X1 $T=1284780 1480510 0 0 $X=1284778 $Y=1480258
X2626 276 12222 283 24 12066 25 12409 AO22X1 $T=1284780 1510030 1 0 $X=1284778 $Y=1506090
X2627 294 11496 285 24 12226 25 12394 AO22X1 $T=1290760 1362430 0 180 $X=1288000 $Y=1358490
X2628 294 11486 285 24 293 25 302 AO22X1 $T=1289840 1355050 1 0 $X=1289838 $Y=1351110
X2629 276 11364 285 24 12392 25 12402 AO22X1 $T=1293060 1443610 1 180 $X=1290300 $Y=1443358
X2630 276 11620 285 24 12463 25 12484 AO22X1 $T=1293060 1480510 0 0 $X=1293058 $Y=1480258
X2631 276 11530 285 24 12350 25 12475 AO22X1 $T=1295820 1414090 1 180 $X=1293060 $Y=1413838
X2632 276 12026 285 24 12408 25 12401 AO22X1 $T=1295820 1436230 0 180 $X=1293060 $Y=1432290
X2633 276 12315 283 24 12379 25 12494 AO22X1 $T=1293520 1510030 1 0 $X=1293518 $Y=1506090
X2634 276 11498 283 24 12470 25 12376 AO22X1 $T=1297660 1399330 0 180 $X=1294900 $Y=1395390
X2635 276 11948 283 24 12483 25 12624 AO22X1 $T=1302260 1510030 1 0 $X=1302258 $Y=1506090
X2636 294 10925 283 24 12578 25 12396 AO22X1 $T=1305020 1369810 1 180 $X=1302260 $Y=1369558
X2637 9934 25 10013 10004 10079 24 10127 NOR4X1 $T=1121940 1458370 0 180 $X=1119640 $Y=1454430
X2638 9993 25 10067 10004 9934 24 10172 NOR4X1 $T=1120560 1458370 0 0 $X=1120558 $Y=1458118
X2639 10179 25 10272 10225 10277 24 103 NOR4X1 $T=1138040 1369810 1 0 $X=1138038 $Y=1365870
X2640 10486 25 10390 10400 10362 24 10466 NOR4X1 $T=1155520 1362430 0 0 $X=1155518 $Y=1362178
X2641 39 25 43 107 44 24 10497 NOR4X1 $T=1159660 1443610 0 180 $X=1157360 $Y=1439670
X2642 10583 25 10511 10505 10614 24 10504 NOR4X1 $T=1173460 1473130 0 0 $X=1173458 $Y=1472878
X2643 181 25 183 88 100 24 11230 NOR4X1 $T=1207040 1524790 0 0 $X=1207038 $Y=1524538
X2644 60 25 12559 74 315 24 10495 NOR4X1 $T=1299960 1399330 0 0 $X=1299958 $Y=1399078
X2645 49 25 24 46 9811 9900 NAND3BX1 $T=1101700 1355050 1 180 $X=1099400 $Y=1354798
X2646 10354 25 24 10289 10187 10279 NAND3BX1 $T=1141720 1473130 1 180 $X=1139420 $Y=1472878
X2647 12500 25 24 10937 275 12364 NAND3BX1 $T=1296280 1391950 0 180 $X=1293980 $Y=1388010
X2648 9738 9674 9687 24 25 XOR2X1 $T=1082840 1414090 1 180 $X=1079620 $Y=1413838
X2649 9679 9738 9754 24 25 XOR2X1 $T=1087900 1377190 0 0 $X=1087898 $Y=1376938
X2650 9827 9813 9809 24 25 XOR2X1 $T=1096180 1362430 0 180 $X=1092960 $Y=1358490
X2651 9811 9829 9821 24 25 XOR2X1 $T=1097560 1369810 0 180 $X=1094340 $Y=1365870
X2652 9831 39 9822 24 25 XOR2X1 $T=1097560 1399330 1 180 $X=1094340 $Y=1399078
X2653 9810 9682 9815 24 25 XOR2X1 $T=1098020 1421470 0 180 $X=1094800 $Y=1417530
X2654 9829 9907 9807 24 25 XOR2X1 $T=1102160 1406710 1 180 $X=1098940 $Y=1406458
X2655 9813 9823 9910 24 25 XOR2X1 $T=1099400 1414090 0 0 $X=1099398 $Y=1413838
X2656 9738 9998 9992 24 25 XOR2X1 $T=1112280 1421470 0 180 $X=1109060 $Y=1417530
X2657 9810 10006 10012 24 25 XOR2X1 $T=1111820 1421470 0 0 $X=1111818 $Y=1421218
X2658 10038 9819 10018 24 25 XOR2X1 $T=1115040 1362430 1 180 $X=1111820 $Y=1362178
X2659 10038 9813 10123 24 25 XOR2X1 $T=1120100 1369810 1 0 $X=1120098 $Y=1365870
X2660 9829 10005 10019 24 25 XOR2X1 $T=1123320 1414090 0 180 $X=1120100 $Y=1410150
X2661 9813 10122 9942 24 25 XOR2X1 $T=1123320 1414090 1 180 $X=1120100 $Y=1413838
X2662 9831 84 9946 24 25 XOR2X1 $T=1124240 1406710 0 180 $X=1121020 $Y=1402770
X2663 9737 77 10179 24 25 XOR2X1 $T=1127000 1377190 1 0 $X=1126998 $Y=1373250
X2664 9762 68 10225 24 25 XOR2X1 $T=1128840 1369810 1 0 $X=1128838 $Y=1365870
X2665 10249 10025 10262 24 25 XOR2X1 $T=1135280 1377190 1 0 $X=1135278 $Y=1373250
X2666 9808 10137 10272 24 25 XOR2X1 $T=1137120 1369810 0 0 $X=1137118 $Y=1369558
X2667 151 10805 10883 24 25 XOR2X1 $T=1180360 1355050 1 0 $X=1180358 $Y=1351110
X2668 11370 11336 11324 24 25 XOR2X1 $T=1216700 1362430 0 180 $X=1213480 $Y=1358490
X2669 11378 199 11394 24 25 XOR2X1 $T=1219000 1362430 1 0 $X=1218998 $Y=1358490
X2670 11479 11391 11432 24 25 XOR2X1 $T=1224060 1369810 0 180 $X=1220840 $Y=1365870
X2671 11450 11448 11490 24 25 XOR2X1 $T=1224520 1377190 0 0 $X=1224518 $Y=1376938
X2672 11543 11684 11699 24 25 XOR2X1 $T=1240160 1428850 0 0 $X=1240158 $Y=1428598
X2673 11581 11787 11807 24 25 XOR2X1 $T=1246600 1362430 1 0 $X=1246598 $Y=1358490
X2674 11737 11795 11890 24 25 XOR2X1 $T=1249360 1458370 0 0 $X=1249358 $Y=1458118
X2675 12117 12077 12067 24 25 XOR2X1 $T=1270520 1399330 1 180 $X=1267300 $Y=1399078
X2676 12185 12199 12086 24 25 XOR2X1 $T=1275120 1465750 1 180 $X=1271900 $Y=1465498
X2677 12230 12203 12216 24 25 XOR2X1 $T=1277880 1399330 1 180 $X=1274660 $Y=1399078
X2678 12250 12184 12072 24 25 XOR2X1 $T=1279720 1458370 0 180 $X=1276500 $Y=1454430
X2679 12241 12346 12341 24 25 XOR2X1 $T=1283400 1399330 1 0 $X=1283398 $Y=1395390
X2680 9815 9687 24 9673 25 9669 OAI21XL $T=1082380 1414090 0 180 $X=1080540 $Y=1410150
X2681 9672 9740 24 9745 25 9668 OAI21XL $T=1083760 1391950 0 0 $X=1083758 $Y=1391698
X2682 10012 9992 24 9673 25 10024 OAI21XL $T=1112740 1421470 1 0 $X=1112738 $Y=1417530
X2683 10003 10029 24 9745 25 10037 OAI21XL $T=1113660 1391950 1 0 $X=1113658 $Y=1388010
X2684 104 10055 24 10164 25 10150 OAI21XL $T=1127920 1399330 1 180 $X=1126080 $Y=1399078
X2685 89 10517 24 10164 25 10464 OAI21XL $T=1164720 1369810 1 180 $X=1162880 $Y=1369558
X2686 10872 10814 24 10875 25 10908 OAI21XL $T=1182660 1377190 1 0 $X=1182658 $Y=1373250
X2687 10935 11077 24 11088 25 173 OAI21XL $T=1197380 1355050 0 0 $X=1197378 $Y=1354798
X2688 11337 11297 24 11328 25 11211 OAI21XL $T=1216240 1369810 1 180 $X=1214400 $Y=1369558
X2689 11304 11339 24 11172 25 11325 OAI21XL $T=1216240 1391950 0 180 $X=1214400 $Y=1388010
X2690 11320 11520 24 11522 25 11592 OAI21XL $T=1235100 1391950 0 180 $X=1233260 $Y=1388010
X2691 11602 11535 24 11593 25 11695 OAI21XL $T=1236940 1473130 0 0 $X=1236938 $Y=1472878
X2692 11673 11737 24 11602 25 11688 OAI21XL $T=1243380 1458370 1 180 $X=1241540 $Y=1458118
X2693 11799 11764 24 11738 25 11441 OAI21XL $T=1245220 1473130 0 180 $X=1243380 $Y=1469190
X2694 12190 12185 24 12176 25 12100 OAI21XL $T=1272820 1480510 0 180 $X=1270980 $Y=1476570
X2695 11626 12189 24 11617 25 11915 OAI21XL $T=1273740 1450990 1 180 $X=1271900 $Y=1450738
X2696 12176 12065 24 12073 25 12183 OAI21XL $T=1273740 1480510 1 180 $X=1271900 $Y=1480258
X2697 12184 12246 24 12235 25 12217 OAI21XL $T=1280180 1465750 0 180 $X=1278340 $Y=1461810
X2698 10760 10752 10662 24 25 10452 MX2X1 $T=1175760 1406710 0 180 $X=1172080 $Y=1402770
X2699 10760 11224 11188 24 25 11072 MX2X1 $T=1208880 1406710 0 180 $X=1205200 $Y=1402770
X2700 10760 11483 11393 24 25 11250 MX2X1 $T=1226360 1414090 1 180 $X=1222680 $Y=1413838
X2701 10952 12233 12315 24 25 12080 MX2X1 $T=1277880 1524790 0 0 $X=1277878 $Y=1524538
X2702 30 9677 9672 24 25 XOR2XL $T=1078700 1391950 0 180 $X=1075480 $Y=1388010
X2703 9679 9737 9689 24 25 XOR2XL $T=1083300 1377190 0 180 $X=1080080 $Y=1373250
X2704 9811 9808 9742 24 25 XOR2XL $T=1094800 1369810 1 180 $X=1091580 $Y=1369558
X2705 9827 9819 9744 24 25 XOR2XL $T=1096180 1362430 1 180 $X=1092960 $Y=1362178
X2706 43 9816 9740 24 25 XOR2XL $T=1097100 1391950 1 180 $X=1093880 $Y=1391698
X2707 46 9810 9820 24 25 XOR2XL $T=1098020 1369810 1 180 $X=1094800 $Y=1369558
X2708 9907 9842 9903 24 25 XOR2XL $T=1102620 1399330 0 180 $X=1099400 $Y=1395390
X2709 46 9762 9922 24 25 XOR2XL $T=1102620 1369810 1 0 $X=1102618 $Y=1365870
X2710 10005 9842 9950 24 25 XOR2XL $T=1111820 1399330 1 180 $X=1108600 $Y=1399078
X2711 59 9677 10003 24 25 XOR2XL $T=1109520 1384570 0 0 $X=1109518 $Y=1384318
X2712 9999 9831 9812 24 25 XOR2XL $T=1112740 1377190 0 180 $X=1109520 $Y=1373250
X2713 9810 68 10021 24 25 XOR2XL $T=1111360 1369810 1 0 $X=1111358 $Y=1365870
X2714 9999 10025 10001 24 25 XOR2XL $T=1114580 1369810 1 180 $X=1111360 $Y=1369558
X2715 60 9816 10029 24 25 XOR2XL $T=1111820 1391950 0 0 $X=1111818 $Y=1391698
X2716 9738 77 10071 24 25 XOR2XL $T=1116880 1377190 1 0 $X=1116878 $Y=1373250
X2717 9829 10137 10145 24 25 XOR2XL $T=1128840 1369810 0 0 $X=1128838 $Y=1369558
X2718 10033 39 98 24 25 XOR2XL $T=1137120 1355050 1 0 $X=1137118 $Y=1351110
X2719 10137 9907 99 24 25 XOR2XL $T=1137120 1355050 0 0 $X=1137118 $Y=1354798
X2720 77 59 10362 24 25 XOR2XL $T=1142640 1369810 1 0 $X=1142638 $Y=1365870
X2721 68 60 10377 24 25 XOR2XL $T=1149080 1362430 0 180 $X=1145860 $Y=1358490
X2722 10137 10005 10390 24 25 XOR2XL $T=1146320 1362430 0 0 $X=1146318 $Y=1362178
X2723 10033 84 10400 24 25 XOR2XL $T=1147240 1369810 1 0 $X=1147238 $Y=1365870
X2724 76 74 10486 24 25 XOR2XL $T=1157820 1362430 0 180 $X=1154600 $Y=1358490
X2725 10742 10732 10728 24 25 XOR2XL $T=1174380 1399330 0 180 $X=1171160 $Y=1395390
X2726 10762 10724 10733 24 25 XOR2XL $T=1175760 1421470 0 180 $X=1172540 $Y=1417530
X2727 10737 10731 10780 24 25 XOR2XL $T=1173920 1428850 1 0 $X=1173918 $Y=1424910
X2728 10798 10779 10752 24 25 XOR2XL $T=1177140 1406710 1 180 $X=1173920 $Y=1406458
X2729 158 10909 10969 24 25 XOR2XL $T=1188640 1436230 1 0 $X=1188638 $Y=1432290
X2730 10887 11042 10946 24 25 XOR2XL $T=1194160 1436230 1 180 $X=1190940 $Y=1435978
X2731 11178 10848 11108 24 25 XOR2XL $T=1205660 1399330 1 180 $X=1202440 $Y=1399078
X2732 11203 11110 11119 24 25 XOR2XL $T=1208880 1450990 0 180 $X=1205660 $Y=1447050
X2733 11227 11246 11199 24 25 XOR2XL $T=1210260 1465750 1 180 $X=1207040 $Y=1465498
X2734 11316 11309 11338 24 25 XOR2XL $T=1213480 1502650 1 0 $X=1213478 $Y=1498710
X2735 11317 11319 11345 24 25 XOR2XL $T=1213480 1524790 1 0 $X=1213478 $Y=1520850
X2736 11313 11301 11224 24 25 XOR2XL $T=1217160 1406710 0 180 $X=1213940 $Y=1402770
X2737 11362 11367 11382 24 25 XOR2XL $T=1217160 1495270 1 0 $X=1217158 $Y=1491330
X2738 11383 11351 11358 24 25 XOR2XL $T=1223140 1473130 0 0 $X=1223138 $Y=1472878
X2739 189 11485 11483 24 25 XOR2XL $T=1226360 1414090 1 0 $X=1226358 $Y=1410150
X2740 11614 11601 11510 24 25 XOR2XL $T=1234180 1517410 0 180 $X=1230960 $Y=1513470
X2741 11690 11666 11597 24 25 XOR2XL $T=1239700 1517410 0 180 $X=1236480 $Y=1513470
X2742 11647 11660 11607 24 25 XOR2XL $T=1237860 1414090 0 0 $X=1237858 $Y=1413838
X2743 11775 11683 11698 24 25 XOR2XL $T=1245220 1406710 0 180 $X=1242000 $Y=1402770
X2744 11739 11760 11742 24 25 XOR2XL $T=1245220 1517410 0 180 $X=1242000 $Y=1513470
X2745 11925 11892 11876 24 25 XOR2XL $T=1254880 1399330 1 180 $X=1251660 $Y=1399078
X2746 11918 11891 11966 24 25 XOR2XL $T=1257640 1510030 0 0 $X=1257638 $Y=1509778
X2747 12053 12019 12035 24 25 XOR2XL $T=1265460 1406710 0 180 $X=1262240 $Y=1402770
X2748 12014 11944 12092 24 25 XOR2XL $T=1265460 1517410 1 0 $X=1265458 $Y=1513470
X2749 12030 12099 12063 24 25 XOR2XL $T=1269140 1517410 1 180 $X=1265920 $Y=1517158
X2750 12173 12105 12200 24 25 XOR2XL $T=1271440 1517410 1 0 $X=1271438 $Y=1513470
X2751 12228 12229 12233 24 25 XOR2XL $T=1280180 1517410 0 180 $X=1276960 $Y=1513470
X2752 10473 10267 25 10492 10505 10511 10465 10454 24 AOI222XL $T=1155060 1487890 1 0 $X=1155058 $Y=1483950
X2753 11907 11249 25 11580 11921 241 11327 11932 24 AOI222XL $T=1252580 1436230 1 0 $X=1252578 $Y=1432290
X2754 12224 11249 25 11580 12172 272 11327 12254 24 AOI222XL $T=1276500 1436230 1 0 $X=1276498 $Y=1432290
X2755 10953 156 10919 24 25 11041 AO21X1 $T=1189100 1362430 0 0 $X=1189098 $Y=1362178
X2756 11016 11085 11027 24 25 10958 AO21X1 $T=1193700 1377190 0 180 $X=1191400 $Y=1373250
X2757 11236 11232 11211 24 25 11085 AO21X1 $T=1209340 1377190 0 180 $X=1207040 $Y=1373250
X2758 11533 11670 11631 24 25 11598 AO21X1 $T=1236940 1391950 1 180 $X=1234640 $Y=1391698
X2759 11249 12212 12220 24 25 12109 AO21X1 $T=1277420 1399330 0 180 $X=1275120 $Y=1395390
X2760 11249 12231 12225 24 25 12112 AO21X1 $T=1278340 1406710 1 180 $X=1276040 $Y=1406458
X2761 9736 9816 25 9810 9739 24 38 AOI22XL $T=1095720 1384570 0 180 $X=1092960 $Y=1380630
X2762 9736 9836 25 9813 9739 24 47 AOI22XL $T=1098020 1384570 0 0 $X=1098018 $Y=1384318
X2763 9736 9842 25 9829 9739 24 9824 AOI22XL $T=1098480 1384570 1 0 $X=1098478 $Y=1380630
X2764 9736 9899 25 9831 9739 24 50 AOI22XL $T=1098940 1391950 1 0 $X=1098938 $Y=1388010
X2765 10899 10798 25 10857 10854 24 10873 AOI22XL $T=1183120 1406710 0 180 $X=1180360 $Y=1402770
X2766 10899 10887 25 10865 10854 24 10886 AOI22XL $T=1183120 1443610 1 180 $X=1180360 $Y=1443358
X2767 10899 10762 25 10884 10854 24 10809 AOI22XL $T=1184040 1414090 1 180 $X=1181280 $Y=1413838
X2768 10899 10742 25 10933 10854 24 10967 AOI22XL $T=1184960 1399330 0 0 $X=1184958 $Y=1399078
X2769 10899 10737 25 10934 10854 24 10968 AOI22XL $T=1184960 1421470 0 0 $X=1184958 $Y=1421218
X2770 166 10615 25 10460 10964 24 10811 AOI22XL $T=1193240 1524790 1 180 $X=1190480 $Y=1524538
X2771 11073 158 25 10949 11098 24 11109 AOI22XL $T=1196920 1436230 0 0 $X=1196918 $Y=1435978
X2772 11073 11203 25 11201 11098 24 11226 AOI22XL $T=1208880 1443610 1 180 $X=1206120 $Y=1443358
X2773 10899 11227 25 11218 11098 24 11228 AOI22XL $T=1208880 1465750 0 180 $X=1206120 $Y=1461810
X2774 10899 11178 25 11247 11249 24 11118 AOI22XL $T=1207960 1399330 0 0 $X=1207958 $Y=1399078
X2775 10899 189 25 11326 11249 24 11225 AOI22XL $T=1213020 1428850 0 0 $X=1213018 $Y=1428598
X2776 10899 11362 25 11330 11098 24 11363 AOI22XL $T=1218080 1487890 1 180 $X=1215320 $Y=1487638
X2777 11327 11313 25 11318 11249 24 11340 AOI22XL $T=1216700 1414090 1 0 $X=1216698 $Y=1410150
X2778 10899 11317 25 11307 11098 24 11398 AOI22XL $T=1217160 1517410 1 0 $X=1217158 $Y=1513470
X2779 11073 11383 25 11315 11098 24 11333 AOI22XL $T=1219000 1473130 1 0 $X=1218998 $Y=1469190
X2780 10899 11316 25 11238 11098 24 11389 AOI22XL $T=1224060 1502650 0 0 $X=1224058 $Y=1502398
X2781 10899 11614 25 11381 11098 24 11603 AOI22XL $T=1235100 1510030 0 180 $X=1232340 $Y=1506090
X2782 10899 11739 25 11693 11098 24 11696 AOI22XL $T=1243380 1502650 1 180 $X=1240620 $Y=1502398
X2783 10899 11690 25 11740 11098 24 11613 AOI22XL $T=1241080 1510030 1 0 $X=1241078 $Y=1506090
X2784 10899 11918 25 11930 11098 24 11901 AOI22XL $T=1253500 1510030 1 0 $X=1253498 $Y=1506090
X2785 10899 12014 25 12023 11098 24 11929 AOI22XL $T=1259480 1510030 1 0 $X=1259478 $Y=1506090
X2786 12017 10899 25 12063 11098 24 12074 AOI22XL $T=1267300 1495270 1 180 $X=1264540 $Y=1495018
X2787 10899 269 25 12215 11098 24 12104 AOI22XL $T=1277880 1510030 0 180 $X=1275120 $Y=1506090
X2788 10899 12228 25 12192 11098 24 12089 AOI22XL $T=1278340 1502650 1 180 $X=1275580 $Y=1502398
X2789 12055 10775 12221 25 12212 24 XOR3X1 $T=1282940 1414090 0 180 $X=1275120 $Y=1410150
X2790 12170 12184 24 25 12168 NAND2BXL $T=1272820 1458370 0 180 $X=1270980 $Y=1454430
X2791 10775 10713 10885 10904 25 24 10884 ADDFXL $T=1176220 1421470 1 0 $X=1176218 $Y=1417530
X2792 10775 10508 10876 10924 25 24 10933 ADDFXL $T=1177600 1414090 1 0 $X=1177598 $Y=1410150
X2793 10775 10761 10888 10920 25 24 10949 ADDFXL $T=1178060 1436230 1 0 $X=1178058 $Y=1432290
X2794 10775 10717 10920 10885 25 24 10934 ADDFXL $T=1178980 1428850 0 0 $X=1178978 $Y=1428598
X2795 10775 10452 10904 10876 25 24 10857 ADDFXL $T=1190020 1406710 1 180 $X=1180820 $Y=1406458
X2796 10936 10807 10910 10888 25 24 10865 ADDFXL $T=1190480 1450990 0 180 $X=1181280 $Y=1447050
X2797 11068 10950 11173 10910 25 24 11201 ADDFXL $T=1196000 1458370 1 0 $X=1195998 $Y=1454430
X2798 11084 11029 11189 11173 25 24 11218 ADDFXL $T=1198300 1473130 0 0 $X=1198298 $Y=1472878
X2799 11128 11076 11207 11229 25 24 11238 ADDFXL $T=1200140 1510030 1 0 $X=1200138 $Y=1506090
X2800 10775 11072 11217 11237 25 24 11318 ADDFXL $T=1201060 1414090 0 0 $X=1201058 $Y=1413838
X2801 11129 11198 11231 11207 25 24 11307 ADDFXL $T=1201980 1524790 1 0 $X=1201978 $Y=1520850
X2802 10775 10944 10924 11217 25 24 11247 ADDFXL $T=1202440 1406710 0 0 $X=1202438 $Y=1406458
X2803 11177 11195 11229 11261 25 24 11330 ADDFXL $T=1202440 1487890 0 0 $X=1202438 $Y=1487638
X2804 11176 11167 11261 11189 25 24 11315 ADDFXL $T=1204740 1480510 1 0 $X=1204738 $Y=1476570
X2805 10775 11250 11237 11462 25 24 11326 ADDFXL $T=1216240 1428850 1 0 $X=1216238 $Y=1424910
X2806 11531 11476 11433 11231 25 24 11381 ADDFXL $T=1228200 1524790 0 180 $X=1219000 $Y=1520850
X2807 11627 11658 11686 11433 25 24 11740 ADDFXL $T=1235100 1524790 1 0 $X=1235098 $Y=1520850
X2808 11642 11532 11700 11686 25 24 11693 ADDFXL $T=1236020 1524790 0 0 $X=1236018 $Y=1524538
X2809 10775 11668 11442 11762 25 24 11935 ADDFXL $T=1236480 1421470 1 0 $X=1236478 $Y=1417530
X2810 10775 11905 11762 11797 25 24 11790 ADDFXL $T=1255800 1414090 1 180 $X=1246600 $Y=1413838
X2811 10775 11873 11797 11926 25 24 11946 ADDFXL $T=1247060 1421470 0 0 $X=1247058 $Y=1421218
X2812 11809 11893 11923 11700 25 24 11930 ADDFXL $T=1248440 1524790 0 0 $X=1248438 $Y=1524538
X2813 11919 11943 12015 11923 25 24 12023 ADDFXL $T=1253960 1532170 1 0 $X=1253958 $Y=1528230
X2814 10775 11957 11926 12049 25 24 12091 ADDFXL $T=1255800 1414090 0 0 $X=1255798 $Y=1413838
X2815 12038 12080 12118 12186 25 24 12192 ADDFXL $T=1264080 1524790 0 0 $X=1264078 $Y=1524538
X2816 12027 12103 12186 12015 25 24 12215 ADDFXL $T=1265920 1532170 0 0 $X=1265918 $Y=1531918
X2817 10775 12181 12049 12221 25 24 12231 ADDFXL $T=1269600 1414090 0 0 $X=1269598 $Y=1413838
X2818 11608 11487 11499 10663 10915 11632 11614 25 24 SDFFRX2 $T=1246600 1487890 1 180 $X=1234180 $Y=1487638
X2819 12109 224 12166 229 10810 270 12241 25 24 SDFFRX2 $T=1267760 1391950 0 0 $X=1267758 $Y=1391698
X2820 12095 11487 12177 11960 10915 12243 12229 25 24 SDFFRX2 $T=1268680 1495270 0 0 $X=1268678 $Y=1495018
X2821 12098 11487 12173 11960 10915 12244 12228 25 24 SDFFRX2 $T=1268680 1502650 1 0 $X=1268678 $Y=1498710
X2822 9673 9671 24 9669 25 9668 9670 OAI211X1 $T=1076860 1399330 1 180 $X=1074560 $Y=1399078
X2823 9673 10014 24 10024 25 10037 10030 OAI211X1 $T=1111820 1399330 1 0 $X=1111818 $Y=1395390
X2824 10587 10801 24 10809 25 10815 10855 OAI211X1 $T=1178060 1414090 0 0 $X=1178058 $Y=1413838
X2825 10050 10801 24 10873 25 10893 10898 OAI211X1 $T=1180820 1399330 1 0 $X=1180818 $Y=1395390
X2826 9924 10801 24 10967 25 11050 11020 OAI211X1 $T=1190940 1399330 0 0 $X=1190938 $Y=1399078
X2827 10032 10801 24 10968 25 11009 11061 OAI211X1 $T=1190940 1421470 0 0 $X=1190938 $Y=1421218
X2828 11023 10801 24 10886 25 11087 11099 OAI211X1 $T=1196000 1443610 1 0 $X=1195998 $Y=1439670
X2829 9997 10801 24 11118 25 11125 11033 OAI211X1 $T=1198300 1399330 1 0 $X=1198298 $Y=1395390
X2830 11062 10801 24 11109 25 11127 11080 OAI211X1 $T=1198300 1428850 0 0 $X=1198298 $Y=1428598
X2831 10796 10801 24 11225 25 11212 11069 OAI211X1 $T=1206580 1428850 0 0 $X=1206578 $Y=1428598
X2832 11255 11321 24 11333 25 11344 11322 OAI211X1 $T=1213480 1473130 1 0 $X=1213478 $Y=1469190
X2833 10632 10801 24 11340 25 11343 11183 OAI211X1 $T=1213940 1399330 0 0 $X=1213938 $Y=1399078
X2834 11213 11321 24 11226 25 11347 11379 OAI211X1 $T=1213940 1443610 0 0 $X=1213938 $Y=1443358
X2835 11104 11321 24 11228 25 11380 11443 OAI211X1 $T=1217160 1465750 1 0 $X=1217158 $Y=1461810
X2836 11223 11321 24 11389 25 11392 11461 OAI211X1 $T=1218540 1502650 1 0 $X=1218538 $Y=1498710
X2837 11197 11321 24 11398 25 11444 11481 OAI211X1 $T=1220380 1510030 0 0 $X=1220378 $Y=1509778
X2838 11171 11321 24 11363 25 11488 11538 OAI211X1 $T=1224060 1487890 0 0 $X=1224058 $Y=1487638
X2839 11585 11321 24 11603 25 11609 11608 OAI211X1 $T=1231880 1487890 0 0 $X=1231878 $Y=1487638
X2840 11596 11321 24 11613 25 11619 11640 OAI211X1 $T=1232800 1495270 0 0 $X=1232798 $Y=1495018
X2841 11685 11321 24 11696 25 11747 11771 OAI211X1 $T=1241080 1495270 0 0 $X=1241078 $Y=1495018
X2842 11886 11321 24 11901 25 11900 11796 OAI211X1 $T=1250280 1502650 1 0 $X=1250278 $Y=1498710
X2843 11321 11888 24 11929 25 11936 12057 OAI211X1 $T=1253500 1487890 0 0 $X=1253498 $Y=1487638
X2844 12062 11321 24 12089 25 12096 12098 OAI211X1 $T=1265920 1502650 1 0 $X=1265918 $Y=1498710
X2845 11222 11321 24 12104 25 12087 12058 OAI211X1 $T=1267300 1502650 0 0 $X=1267298 $Y=1502398
X2846 12012 11321 24 12074 25 12094 12095 OAI211X1 $T=1270060 1495270 0 180 $X=1267760 $Y=1491330
X2847 214 11252 10954 25 11371 11595 24 AOI2BB2X1 $T=1235560 1377190 1 180 $X=1232800 $Y=1376938
X2848 11897 10801 11249 25 11790 11793 24 AOI2BB2X1 $T=1251660 1406710 1 180 $X=1248900 $Y=1406458
X2849 11958 10801 11249 25 11935 11768 24 AOI2BB2X1 $T=1259020 1421470 0 180 $X=1256260 $Y=1417530
X2850 250 11252 10954 25 11875 11961 24 AOI2BB2X1 $T=1261320 1377190 1 180 $X=1258560 $Y=1376938
X2851 12085 10801 11249 25 11946 12059 24 AOI2BB2X1 $T=1267760 1421470 0 180 $X=1265000 $Y=1417530
X2852 260 11252 10954 25 11667 12083 24 AOI2BB2X1 $T=1270060 1377190 1 180 $X=1267300 $Y=1376938
X2853 12204 10801 11249 25 12091 12048 24 AOI2BB2X1 $T=1270060 1406710 1 180 $X=1267300 $Y=1406458
X2854 10033 9831 10129 25 24 XNOR2X1 $T=1125160 1377190 0 180 $X=1121940 $Y=1373250
X2855 10734 146 10759 25 24 XNOR2X1 $T=1173460 1362430 1 0 $X=1173458 $Y=1358490
X2856 10958 10917 10927 25 24 XNOR2X1 $T=1188180 1369810 1 180 $X=1184960 $Y=1369558
X2857 11085 11097 11116 25 24 XNOR2X1 $T=1197840 1377190 1 0 $X=1197838 $Y=1373250
X2858 11041 11169 11175 25 24 XNOR2X1 $T=1200600 1362430 0 0 $X=1200598 $Y=1362178
X2859 11598 11537 11578 25 24 XNOR2X1 $T=1234180 1384570 1 180 $X=1230960 $Y=1384318
X2860 11679 11644 11594 25 24 XNOR2X1 $T=1239700 1377190 0 180 $X=1236480 $Y=1373250
X2861 11688 11639 11669 25 24 XNOR2X1 $T=1241540 1450990 1 180 $X=1238320 $Y=1450738
X2862 11770 11657 11677 25 24 XNOR2X1 $T=1242460 1443610 1 180 $X=1239240 $Y=1443358
X2863 11682 11748 11641 25 24 XNOR2X1 $T=1242460 1369810 1 0 $X=1242458 $Y=1365870
X2864 11670 11734 11749 25 24 XNOR2X1 $T=1242920 1399330 1 0 $X=1242918 $Y=1395390
X2865 11885 11884 11802 25 24 XNOR2X1 $T=1251660 1465750 0 180 $X=1248440 $Y=1461810
X2866 11950 11962 11967 25 24 XNOR2X1 $T=1258100 1458370 0 0 $X=1258098 $Y=1458118
X2867 12100 12088 12070 25 24 XNOR2X1 $T=1268680 1480510 0 180 $X=1265460 $Y=1476570
X2868 9993 25 10067 24 10034 10131 NOR3X1 $T=1123780 1465750 1 180 $X=1121940 $Y=1465498
X2869 10369 25 10488 24 10280 10487 NOR3X1 $T=1156900 1465750 0 180 $X=1155060 $Y=1461810
X2870 10568 25 10474 24 10488 10344 NOR3X1 $T=1159200 1465750 1 180 $X=1157360 $Y=1465498
X2871 10583 25 10511 24 10614 10961 NOR3X1 $T=1190020 1495270 0 0 $X=1190018 $Y=1495018
X2872 166 25 170 24 65 11959 NOR3X1 $T=1261780 1517410 0 0 $X=1261778 $Y=1517158
X2873 10159 10143 10131 24 10127 25 10125 AND4X1 $T=1124700 1465750 0 180 $X=1121940 $Y=1461810
X2874 10868 10866 10947 24 10754 25 10955 AND4X1 $T=1186800 1510030 0 0 $X=1186798 $Y=1509778
X2875 10955 10867 10773 24 10811 25 10931 AND4X1 $T=1189100 1517410 0 0 $X=1189098 $Y=1517158
X2876 11117 11252 11220 24 11233 25 10854 AND4X1 $T=1210720 1450990 1 180 $X=1207960 $Y=1450738
X2877 12046 12012 95 24 11959 25 11302 AND4X1 $T=1260860 1502650 1 180 $X=1258100 $Y=1502398
X2878 10614 10505 10164 24 25 10595 AO21XL $T=1164260 1465750 1 180 $X=1161960 $Y=1465498
X2879 11933 11885 11940 24 25 11950 AO21XL $T=1255340 1465750 1 0 $X=1255338 $Y=1461810
X2880 10183 10188 25 10224 24 10187 AOI21X1 $T=1129300 1480510 0 0 $X=1129298 $Y=1480258
X2881 10274 10267 25 10261 24 10260 AOI21X1 $T=1138960 1480510 1 180 $X=1136660 $Y=1480258
X2882 11388 11232 25 11489 24 11479 AOI21X1 $T=1224980 1377190 1 0 $X=1224978 $Y=1373250
X2883 11513 11582 25 11592 24 11339 AOI21X1 $T=1231420 1399330 0 0 $X=1231418 $Y=1399078
X2884 207 11445 25 11600 24 11581 AOI21X1 $T=1231880 1355050 0 0 $X=1231878 $Y=1354798
X2885 11691 11682 25 11741 24 11679 AOI21X1 $T=1241540 1377190 0 0 $X=1241538 $Y=1376938
X2886 11689 11756 25 11695 24 11738 AOI21X1 $T=1244760 1473130 1 180 $X=1242460 $Y=1472878
X2887 11808 11885 25 11756 24 11737 AOI21X1 $T=1251200 1465750 1 180 $X=1248900 $Y=1465498
X2888 170 10615 25 10964 10882 24 10867 AOI22X1 $T=1191860 1517410 0 180 $X=1189100 $Y=1513470
X2889 174 10615 25 10614 10964 24 10866 AOI22X1 $T=1198760 1510030 0 180 $X=1196000 $Y=1506090
X2890 183 10615 25 10511 10964 24 10773 AOI22X1 $T=1199220 1517410 1 180 $X=1196460 $Y=1517158
X2891 181 10615 25 10583 10964 24 10868 AOI22X1 $T=1201060 1524790 1 180 $X=1198300 $Y=1524538
X2892 11249 11375 25 11368 87 24 11376 AOI22X1 $T=1219460 1436230 0 180 $X=1216700 $Y=1432290
X2893 11800 10899 25 11507 10954 24 11774 AOI22X1 $T=1245680 1391950 1 180 $X=1242920 $Y=1391698
X2894 10396 10760 24 11073 25 NAND2BX1 $T=1196920 1465750 0 0 $X=1196918 $Y=1465498
X2895 11431 11252 24 11523 25 NAND2BX1 $T=1225900 1458370 1 0 $X=1225898 $Y=1454430
X2896 11678 11653 24 11748 25 NAND2BX1 $T=1242920 1369810 0 0 $X=1242918 $Y=1369558
X2897 77 10264 101 24 25 10121 OA21XL $T=1138040 1362430 1 0 $X=1138038 $Y=1358490
X2898 10494 10499 119 24 25 121 OA21XL $T=1156440 1355050 0 0 $X=1156438 $Y=1354798
X2899 10494 10065 119 24 25 128 OA21XL $T=1161500 1355050 0 0 $X=1161498 $Y=1354798
X2900 11184 10817 11196 24 25 10599 OA21XL $T=1208880 1495270 0 180 $X=1206580 $Y=1491330
X2901 195 11336 196 24 25 11378 OA21XL $T=1215780 1355050 0 0 $X=1215778 $Y=1354798
X2902 11502 11543 11649 24 25 11763 OA21XL $T=1242460 1436230 0 0 $X=1242458 $Y=1435978
X2903 9899 39 9671 24 25 XNOR2XL $T=1096180 1399330 0 180 $X=1092960 $Y=1395390
X2904 9836 44 9814 24 25 XNOR2XL $T=1098020 1406710 0 180 $X=1094800 $Y=1402770
X2905 34 9907 54 24 25 XNOR2XL $T=1107220 1355050 1 180 $X=1104000 $Y=1354798
X2906 9836 74 10023 24 25 XNOR2XL $T=1120100 1406710 0 0 $X=1120098 $Y=1406458
X2907 9899 84 10014 24 25 XNOR2XL $T=1123320 1399330 0 180 $X=1120100 $Y=1395390
X2908 34 10005 10120 24 25 XNOR2XL $T=1121940 1355050 0 0 $X=1121938 $Y=1354798
X2909 10892 10817 10874 24 25 XNOR2XL $T=1184040 1495270 0 180 $X=1180820 $Y=1491330
X2910 11445 11525 11586 24 25 XNOR2XL $T=1230500 1355050 1 0 $X=1230498 $Y=1351110
X2911 24 31 45 9900 53 9926 25 OAI31XL $T=1103080 1355050 1 0 $X=1103078 $Y=1351110
X2912 24 10267 10389 10386 10380 10261 25 OAI31XL $T=1148620 1487890 1 180 $X=1146320 $Y=1487638
X2913 24 10520 10457 10475 10471 10226 25 OAI31XL $T=1154140 1450990 1 180 $X=1151840 $Y=1450738
X2914 24 101 11499 11021 11018 11541 25 OAI31XL $T=1226360 1458370 0 0 $X=1226358 $Y=1458118
X2915 10775 11449 11462 11442 24 25 11375 CMPR32X2 $T=1231420 1421470 1 180 $X=1221760 $Y=1421218
X2916 11327 11233 24 11251 25 11354 NAND3BXL $T=1214400 1450990 1 0 $X=1214398 $Y=1447050
X2917 11251 11220 11184 25 24 11431 AOI2BB1X1 $T=1213940 1458370 1 0 $X=1213938 $Y=1454430
X2918 10663 10241 11080 175 10915 158 24 25 SDFFRHQX8 $T=1195080 1436230 1 0 $X=1195078 $Y=1432290
X2919 10663 11028 11322 197 10915 11383 24 25 SDFFRHQX8 $T=1212100 1465750 0 0 $X=1212098 $Y=1465498
X2920 10460 10447 10243 10457 25 10013 24 NAND4BBXL $T=1152760 1458370 1 180 $X=1149540 $Y=1458118
X2921 10882 10505 10961 10960 25 10460 24 NAND4BBXL $T=1188640 1502650 0 0 $X=1188638 $Y=1502398
X2922 174 11230 11222 11215 25 165 24 NAND4BBXL $T=1208880 1517410 0 180 $X=1205660 $Y=1513470
X2923 10854 11098 24 25 BUFX2 $T=1203360 1436230 0 0 $X=1203358 $Y=1435978
X2924 9804 24 10001 9922 9908 55 25 NAND4XL $T=1107220 1362430 1 180 $X=1104920 $Y=1362178
X2925 10463 24 10371 10373 10473 10339 25 NAND4XL $T=1150920 1473130 0 0 $X=1150918 $Y=1472878
X2926 10473 24 10502 10371 10511 10359 25 NAND4XL $T=1156440 1473130 0 0 $X=1156438 $Y=1472878
X2927 10267 24 10505 10460 10490 10380 25 NAND4XL $T=1156440 1495270 1 0 $X=1156438 $Y=1491330
X2928 101 24 10504 10460 10371 11018 25 NAND4XL $T=1192320 1458370 1 180 $X=1190020 $Y=1458118
X2929 10868 24 10866 11070 10773 11117 25 NAND4XL $T=1200600 1510030 1 180 $X=1198300 $Y=1509778
X2930 10241 11043 11022 9741 10810 10918 24 25 10911 SDFFSXL $T=1194620 1480510 0 180 $X=1184040 $Y=1476570
X2931 11028 11204 11106 10663 10810 10959 24 25 11043 SDFFSXL $T=1207040 1480510 1 180 $X=1196460 $Y=1480258
X2932 10952 10962 11022 25 24 193157 TLATX1 $T=1188640 1480510 0 0 $X=1188638 $Y=1480258
X2933 10952 11059 11106 25 24 193158 TLATX1 $T=1195540 1487890 0 0 $X=1195538 $Y=1487638
X2934 11069 10241 10366 10663 10810 193159 189 25 24 SDFFRX4 $T=1195540 1428850 1 0 $X=1195538 $Y=1424910
X2935 10117 24 9920 10046 10126 10141 25 OAI22XL $T=1121020 1391950 0 0 $X=1121018 $Y=1391698
X2936 10185 24 92 10002 89 10113 25 OAI22XL $T=1129300 1377190 1 180 $X=1127000 $Y=1376938
X2937 10238 24 10226 10056 10126 10151 25 OAI22XL $T=1131600 1421470 1 180 $X=1129300 $Y=1421218
X2938 10287 24 10226 10222 10126 10276 25 OAI22XL $T=1139880 1421470 1 180 $X=1137580 $Y=1421218
X2939 10265 24 92 10239 10126 10286 25 OAI22XL $T=1138040 1391950 0 0 $X=1138038 $Y=1391698
X2940 10273 24 9920 10170 104 10257 25 OAI22XL $T=1142180 1399330 0 180 $X=1139880 $Y=1395390
X2941 10340 24 10282 10361 104 10379 25 OAI22XL $T=1143560 1428850 0 0 $X=1143558 $Y=1428598
X2942 10485 24 10226 10446 10126 10519 25 OAI22XL $T=1155060 1436230 1 0 $X=1155058 $Y=1432290
X2943 10960 24 10874 10970 10959 11059 25 OAI22XL $T=1189560 1487890 0 0 $X=1189558 $Y=1487638
X2944 10371 10504 24 10460 25 11021 AND3XL $T=1185420 1465750 0 0 $X=1185418 $Y=1465498
X2945 10460 10937 24 10504 25 10903 AND3XL $T=1187720 1473130 0 180 $X=1185420 $Y=1469190
X2946 10903 24 10371 25 10795 10880 NAND3XL $T=1183120 1480510 0 180 $X=1181280 $Y=1476570
X2947 141 10485 24 10862 10629 10817 25 10781 OAI32X1 $T=1182660 1450990 1 180 $X=1179440 $Y=1450738
X2948 144 10772 142 24 10734 25 OAI2BB1X1 $T=1176680 1355050 1 180 $X=1174380 $Y=1354798
X2949 10180 25 10369 24 74 10348 NOR3XL $T=1146780 1473130 0 180 $X=1144940 $Y=1469190
X2950 10492 25 10511 24 10583 10490 NOR3XL $T=1161960 1487890 1 180 $X=1160120 $Y=1487638
X2951 10624 25 10371 24 10460 10455 NOR3XL $T=1164720 1473130 0 180 $X=1162880 $Y=1469190
X2952 10267 25 10505 24 10624 10795 NOR3XL $T=1172540 1480510 1 0 $X=1172538 $Y=1476570
X2953 9736 9677 9738 9739 24 25 33 AO22XL $T=1081920 1384570 0 0 $X=1081918 $Y=1384318
X2954 9830 9995 65 9805 24 25 10075 AO22XL $T=1109980 1495270 1 0 $X=1109978 $Y=1491330
X2955 9830 10169 88 9805 24 25 10017 AO22XL $T=1128380 1510030 0 180 $X=1125620 $Y=1506090
X2956 9830 10280 100 9805 24 25 10189 AO22XL $T=1140340 1495270 1 180 $X=1137580 $Y=1495018
X2957 10387 10343 111 9805 24 25 10347 AO22XL $T=1149080 1517410 1 180 $X=1146320 $Y=1517158
X2958 9830 10596 124 10578 24 25 10626 AO22XL $T=1161500 1495270 0 0 $X=1161498 $Y=1495018
X2959 10578 133 9998 10387 24 25 10536 AO22XL $T=1166100 1532170 0 180 $X=1163340 $Y=1528230
X2960 10578 145 10122 10387 24 25 10634 AO22XL $T=1174840 1532170 0 180 $X=1172080 $Y=1528230
X2961 10187 24 10287 25 10146 10340 NAND3X1 $T=1139880 1428850 0 0 $X=1139878 $Y=1428598
X2962 10492 24 10467 25 10373 10624 NAND3X1 $T=1163800 1480510 1 0 $X=1163798 $Y=1476570
X2963 44 25 10005 30 10281 24 10247 NOR4XL $T=1141260 1443610 0 180 $X=1138960 $Y=1439670
X2964 10371 25 10343 10180 10447 24 10169 NOR4XL $T=1150460 1465750 1 180 $X=1148160 $Y=1465498
X2965 10568 25 10474 127 10496 24 84 NOR4XL $T=1161960 1458370 1 0 $X=1161958 $Y=1454430
X2966 9898 24 9821 9809 9908 51 25 NAND4X1 $T=1099400 1362430 0 0 $X=1099398 $Y=1362178
X2967 81 24 10120 83 85 10178 25 NAND4X1 $T=1121020 1355050 1 0 $X=1121018 $Y=1351110
X2968 10129 24 10123 51 10121 10182 25 NAND4X1 $T=1123320 1362430 1 180 $X=1121020 $Y=1362178
X2969 10262 24 10018 55 10121 10277 25 NAND4X1 $T=1137580 1362430 0 0 $X=1137578 $Y=1362178
X2970 10353 24 10338 10186 10238 10282 25 NAND4X1 $T=1142180 1450990 1 180 $X=1139880 $Y=1450738
X2971 10359 24 10339 10260 10251 10255 25 NAND4X1 $T=1142180 1473130 0 180 $X=1139880 $Y=1469190
X2972 10125 24 10281 10344 10348 10266 25 NAND4X1 $T=1140800 1465750 1 0 $X=1140798 $Y=1461810
X2973 10454 24 10374 10373 10266 10354 25 NAND4X1 $T=1147240 1473130 1 180 $X=1144940 $Y=1472878
X2974 10497 24 10495 10496 10487 10475 25 NAND4X1 $T=1157360 1450990 0 180 $X=1155060 $Y=1447050
X2975 10172 24 10504 10501 10271 10520 25 NAND4X1 $T=1156440 1458370 0 0 $X=1156438 $Y=1458118
X2976 10389 10386 25 10467 10371 24 10374 AOI2BB2XL $T=1153220 1480510 0 180 $X=1150460 $Y=1476570
X2977 10178 10377 25 110 10065 10376 24 NOR4BX1 $T=1148160 1355050 1 180 $X=1144940 $Y=1354798
X2978 9742 9689 9744 24 25 9804 AND3X2 $T=1085140 1369810 1 0 $X=1085138 $Y=1365870
X2979 9812 9754 9820 24 25 9898 AND3X2 $T=1094340 1377190 1 0 $X=1094338 $Y=1373250
X2980 10180 10260 10159 24 25 10289 AND3X2 $T=1138500 1480510 1 0 $X=1138498 $Y=1476570
X2981 10230 25 10266 10270 24 10254 10227 AOI211X1 $T=1139880 1465750 1 180 $X=1137580 $Y=1465498
X2982 10275 10243 24 10271 10268 10263 25 NAND4BX1 $T=1139880 1487890 1 180 $X=1137120 $Y=1487638
X2983 60 59 84 25 24 10247 OR3XL $T=1132520 1443610 1 0 $X=1132518 $Y=1439670
X2984 76 10033 10137 68 25 24 10264 OR4X1 $T=1129300 1362430 1 0 $X=1129298 $Y=1358490
X2985 9807 9687 9815 25 24 9840 OR3X2 $T=1093420 1414090 0 0 $X=1093418 $Y=1413838
X2986 10019 9992 10012 25 24 9996 OR3X2 $T=1114120 1414090 1 180 $X=1111360 $Y=1413838
X2987 39 43 9907 25 24 10079 OR3X2 $T=1112280 1450990 1 0 $X=1112278 $Y=1447050
X2988 10071 10021 10145 25 24 10157 OR3X2 $T=1122860 1369810 0 0 $X=1122858 $Y=1369558
X2989 9673 25 9910 9933 24 9839 9927 AOI211XL $T=1107220 1406710 1 180 $X=1104920 $Y=1406458
X2990 9673 25 9942 9933 24 10022 10031 AOI211XL $T=1111820 1406710 0 0 $X=1111818 $Y=1406458
X2991 9903 9745 25 9822 9673 24 9670 9932 AOI221XL $T=1102620 1399330 0 0 $X=1102618 $Y=1399078
X2992 9950 9745 25 9946 9673 24 10030 10039 AOI221XL $T=1111820 1399330 0 0 $X=1111818 $Y=1399078
X2993 10006 24 25 60 BUFX4 $T=1112280 1436230 0 180 $X=1109980 $Y=1432290
X2994 9998 24 25 59 BUFX4 $T=1110900 1443610 1 0 $X=1110898 $Y=1439670
X2995 9996 9946 9942 24 9910 9822 9840 25 9939 OAI33X1 $T=1108600 1414090 0 180 $X=1104920 $Y=1410150
X2996 34 41 9824 24 25 37 OAI2BB1XL $T=1097100 1355050 0 180 $X=1094800 $Y=1351110
X2997 9674 24 30 25 CLKBUFX8 $T=1092960 1421470 0 0 $X=1092958 $Y=1421218
.ENDS
***************************************
.SUBCKT ICV_31 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18
** N=18 EP=18 IP=21 FDC=0
X0 1 2 3 4 5 6 7 8 9 10 SDFFNSRXL $T=-11960 0 0 0 $X=-11962 $Y=-252
X1 11 12 13 14 15 16 8 17 9 MXI4X1 $T=0 0 0 0 $X=-2 $Y=-252
.ENDS
***************************************
.SUBCKT ICV_32 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18
** N=18 EP=18 IP=21 FDC=0
X0 1 2 3 4 5 6 7 8 9 10 SDFFNSRXL $T=0 0 0 0 $X=-2 $Y=-252
X1 11 12 13 14 15 16 8 17 9 MXI4X1 $T=11960 0 0 0 $X=11958 $Y=-252
.ENDS
***************************************
.SUBCKT CLKINVX16 A VSS VDD Y
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI21XL A1 VDD A0 B0 VSS Y
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INVX16 A Y VSS VDD
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI32XL A2 A1 VDD A0 B0 B1 VSS Y
** N=9 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI32X1 A2 A1 VDD A0 B0 B1 VSS Y
** N=9 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI2BB1XL A0N A1N VDD B0 Y VSS
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI221X1 B1 B0 VSS A0 A1 VDD C0 Y
** N=9 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR2XL A B VSS VDD Y
** N=6 EP=5 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI221X2 B0 B1 VSS A0 A1 C0 Y VDD
** N=9 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI32XL A2 A1 VSS A0 B0 Y VDD B1
** N=9 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MX3XL S0 B A S1 C VSS VDD Y
** N=9 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MXI3X1 A S0 B C VSS VDD S1 Y
** N=9 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MXI2XL B S0 Y A VSS VDD
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUFX16 A Y VDD VSS
** N=5 EP=4 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MXI3XL A S0 B C VSS VDD S1 Y
** N=9 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI221X4 B1 B0 A0 A1 C0 Y VSS VDD
** N=9 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OA22XL A1 A0 B0 B1 VSS VDD Y
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MX3X1 C S0 B A S1 VSS VDD Y
** N=9 EP=8 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI21X1 A1 A0 VSS B0 VDD Y
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI211XL A1 VSS A0 C0 VDD B0 Y
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR3BXL AN C VDD B VSS Y
** N=7 EP=6 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI222XL B1 B0 VSS A0 A1 VDD C1 C0 Y
** N=10 EP=9 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI31X1 A2 A1 VDD A0 B0 VSS Y
** N=8 EP=7 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_33 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42 43 44
+ 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64
+ 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84
+ 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104
+ 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124
+ 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144
+ 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164
+ 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184
+ 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204
+ 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223 224
+ 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242 243 244
+ 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261 262 263 264
+ 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281 282 283 284
+ 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300 301 302 303 304
+ 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321 322 323 324
+ 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341 342 343 344
+ 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361 362 363 364
+ 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381 382 383 384
+ 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401 402 403 404
+ 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421 422 423 424
+ 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441 442 443 444
+ 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461 462 463 464
+ 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480 481 482 483 484
+ 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500 501 502 503 504
+ 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520 521 522 523 524
+ 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540 541 542 543 544
+ 545 546 547 548 549 550 551 552 553 554 555 556 557 558 559 560 561 562 563 564
+ 565 566 567 568 569 570 571 572 573 574 575 576 577 578 579 580 581 582 583 584
+ 585 586 587 588 589 590 591 592 593 594 595 596 597 598 599 600 601 602 603 604
+ 605 606 607 608 609 610 611 612 613 614 615 616 617 618 619 620 621 622 623 624
+ 625 626 627 628 629 630 631 632 633 634 635 636 637 638 639 640 641 642 643 644
+ 645 3920
** N=173261 EP=622 IP=35759 FDC=0
X0 8916 8864 25 26 8860 OR2X1 $T=1060760 1185310 0 180 $X=1058920 $Y=1181370
X1 8748 8885 25 26 8863 OR2X1 $T=1060760 1074610 0 0 $X=1060758 $Y=1074358
X2 8827 8885 25 26 9130 OR2X1 $T=1087440 1074610 1 0 $X=1087438 $Y=1070670
X3 8732 9509 25 26 9277 OR2X1 $T=1104000 1185310 1 180 $X=1102160 $Y=1185058
X4 9773 9737 25 26 9826 OR2X1 $T=1114580 1222210 0 0 $X=1114578 $Y=1221958
X5 98 9871 25 26 10139 OR2X1 $T=1131600 1296010 0 0 $X=1131598 $Y=1295758
X6 11164 11139 25 26 11074 OR2X1 $T=1183120 1340290 0 180 $X=1181280 $Y=1336350
X7 10850 220 25 26 222 OR2X1 $T=1229580 1347670 1 0 $X=1229578 $Y=1343730
X8 277 11626 25 26 13026 OR2X1 $T=1271900 1325530 1 0 $X=1271898 $Y=1321590
X9 13389 13361 25 26 13478 OR2X1 $T=1289840 1096750 1 0 $X=1289838 $Y=1092810
X10 26 25 9519 TIELO $T=1101700 1310770 0 0 $X=1101698 $Y=1310518
X11 26 25 13518 TIEHI $T=1330320 1303390 0 0 $X=1330318 $Y=1303138
X12 26 25 13391 TIEHI $T=1355620 1332910 0 0 $X=1355618 $Y=1332658
X13 26 25 13901 TIEHI $T=1358380 1104130 0 0 $X=1358378 $Y=1103878
X14 26 25 13354 TIEHI $T=1368040 1177930 0 0 $X=1368038 $Y=1177678
X15 26 25 13441 TIEHI $T=1368960 1281250 1 0 $X=1368958 $Y=1277310
X16 26 25 13374 TIEHI $T=1374480 1170550 1 0 $X=1374478 $Y=1166610
X17 26 25 13746 TIEHI $T=1381840 1244350 1 0 $X=1381838 $Y=1240410
X18 26 25 13694 TIEHI $T=1384600 1155790 1 0 $X=1384598 $Y=1151850
X19 26 25 13690 TIEHI $T=1385060 1185310 0 0 $X=1385058 $Y=1185058
X20 26 25 13534 TIEHI $T=1389200 1266490 0 0 $X=1389198 $Y=1266238
X21 26 25 13738 TIEHI $T=1389660 1207450 0 0 $X=1389658 $Y=1207198
X22 26 25 13660 TIEHI $T=1390580 1251730 0 0 $X=1390578 $Y=1251478
X23 26 25 13671 TIEHI $T=1392420 1141030 1 0 $X=1392418 $Y=1137090
X24 26 25 13712 TIEHI $T=1397940 1192690 0 0 $X=1397938 $Y=1192438
X25 26 25 13736 TIEHI $T=1400240 1296010 1 0 $X=1400238 $Y=1292070
X26 26 25 13677 TIEHI $T=1401160 1118890 0 0 $X=1401158 $Y=1118638
X27 26 25 13744 TIEHI $T=1401620 1229590 1 0 $X=1401618 $Y=1225650
X28 26 25 13734 TIEHI $T=1403460 1126270 0 0 $X=1403458 $Y=1126018
X29 26 25 13741 TIEHI $T=1405300 1332910 1 0 $X=1405298 $Y=1328970
X30 26 25 13707 TIEHI $T=1407600 1259110 1 0 $X=1407598 $Y=1255170
X31 26 25 13745 TIEHI $T=1408060 1229590 0 0 $X=1408058 $Y=1229338
X32 26 25 13735 TIEHI $T=1408520 1163170 0 0 $X=1408518 $Y=1162918
X33 26 25 13890 TIEHI $T=1411740 1347670 1 0 $X=1411738 $Y=1343730
X34 26 25 13892 TIEHI $T=1419100 1207450 1 0 $X=1419098 $Y=1203510
X35 26 25 13875 TIEHI $T=1420020 1222210 1 0 $X=1420018 $Y=1218270
X36 26 25 13906 TIEHI $T=1423700 1126270 0 0 $X=1423698 $Y=1126018
X37 26 25 13924 TIEHI $T=1427380 1318150 0 0 $X=1427378 $Y=1317898
X38 26 25 14022 TIEHI $T=1428300 1155790 1 0 $X=1428298 $Y=1151850
X39 26 25 13948 TIEHI $T=1429680 1251730 1 0 $X=1429678 $Y=1247790
X40 26 25 14403 TIEHI $T=1431980 1111510 1 0 $X=1431978 $Y=1107570
X41 26 25 14136 TIEHI $T=1431980 1133650 0 0 $X=1431978 $Y=1133398
X42 26 25 14233 TIEHI $T=1446240 1310770 0 0 $X=1446238 $Y=1310518
X43 26 25 14149 TIEHI $T=1448080 1288630 1 0 $X=1448078 $Y=1284690
X44 26 25 14270 TIEHI $T=1449920 1141030 1 0 $X=1449918 $Y=1137090
X45 26 25 14195 TIEHI $T=1454060 1303390 1 0 $X=1454058 $Y=1299450
X46 26 25 14391 TIEHI $T=1460500 1332910 1 0 $X=1460498 $Y=1328970
X47 26 25 14502 TIEHI $T=1461880 1296010 1 0 $X=1461878 $Y=1292070
X48 26 25 14496 TIEHI $T=1469700 1229590 0 0 $X=1469698 $Y=1229338
X49 26 25 14546 TIEHI $T=1469700 1325530 1 0 $X=1469698 $Y=1321590
X50 26 25 14405 TIEHI $T=1470160 1236970 0 0 $X=1470158 $Y=1236718
X51 26 25 14466 TIEHI $T=1470620 1273870 0 0 $X=1470618 $Y=1273618
X52 26 25 14663 TIEHI $T=1473840 1155790 1 0 $X=1473838 $Y=1151850
X53 26 25 14544 TIEHI $T=1474300 1192690 0 0 $X=1474298 $Y=1192438
X54 26 25 444 TIEHI $T=1475680 1347670 1 0 $X=1475678 $Y=1343730
X55 26 25 14586 TIEHI $T=1480740 1177930 0 0 $X=1480738 $Y=1177678
X56 26 25 14671 TIEHI $T=1482580 1303390 0 0 $X=1482578 $Y=1303138
X57 26 25 14691 TIEHI $T=1483500 1200070 0 0 $X=1483498 $Y=1199818
X58 26 25 14580 TIEHI $T=1483500 1259110 0 0 $X=1483498 $Y=1258858
X59 26 25 14581 TIEHI $T=1483500 1281250 0 0 $X=1483498 $Y=1280998
X60 26 25 14838 TIEHI $T=1483960 1229590 1 0 $X=1483958 $Y=1225650
X61 26 25 14623 TIEHI $T=1484420 1185310 0 0 $X=1484418 $Y=1185058
X62 26 25 14839 TIEHI $T=1484880 1163170 0 0 $X=1484878 $Y=1162918
X63 26 25 14731 TIEHI $T=1487180 1207450 0 0 $X=1487178 $Y=1207198
X64 26 25 14801 TIEHI $T=1488560 1266490 1 0 $X=1488558 $Y=1262550
X65 26 25 15035 TIEHI $T=1496380 1340290 1 0 $X=1496378 $Y=1336350
X66 9681 9375 26 25 9510 NOR2BX1 $T=1110440 1244350 1 180 $X=1108600 $Y=1244098
X67 10287 10207 26 25 10042 NOR2BX1 $T=1135280 1089370 0 180 $X=1133440 $Y=1085430
X68 10222 10299 26 25 10192 NOR2BX1 $T=1135740 1104130 1 180 $X=1133900 $Y=1103878
X69 10192 10207 26 25 10230 NOR2BX1 $T=1134360 1111510 1 0 $X=1134358 $Y=1107570
X70 10255 10299 26 25 10287 NOR2BX1 $T=1139420 1089370 1 0 $X=1139418 $Y=1085430
X71 10398 10207 26 25 10406 NOR2BX1 $T=1144020 1089370 1 0 $X=1144018 $Y=1085430
X72 10288 10207 26 25 10438 NOR2BX1 $T=1144940 1118890 0 0 $X=1144938 $Y=1118638
X73 11211 11074 26 25 158 NOR2BX1 $T=1184040 1347670 1 180 $X=1182200 $Y=1347418
X74 11464 11030 26 25 11404 NOR2BX1 $T=1198300 1081990 0 180 $X=1196460 $Y=1078050
X75 11566 10951 26 25 11464 NOR2BX1 $T=1205200 1081990 1 0 $X=1205198 $Y=1078050
X76 11627 10605 26 25 11596 NOR2BX1 $T=1208880 1089370 0 180 $X=1207040 $Y=1085430
X77 11838 10951 26 25 11738 NOR2BX1 $T=1215320 1059850 1 180 $X=1213480 $Y=1059598
X78 11738 11030 26 25 11808 NOR2BX1 $T=1213940 1059850 1 0 $X=1213938 $Y=1055910
X79 11958 11030 26 25 12002 NOR2BX1 $T=1223140 1045090 1 0 $X=1223138 $Y=1041150
X80 458 560 26 25 16027 NOR2BX1 $T=1529960 1347670 0 0 $X=1529958 $Y=1347418
X81 15982 369 26 25 15949 NOR2BX1 $T=1532260 1200070 0 180 $X=1530420 $Y=1196130
X82 398 16076 26 25 16088 NOR2BX1 $T=1540080 1310770 1 180 $X=1538240 $Y=1310518
X83 546 16076 26 25 16008 NOR2BX1 $T=1540080 1318150 0 180 $X=1538240 $Y=1314210
X84 536 16092 26 25 16164 NOR2BX1 $T=1541920 1177930 0 0 $X=1541918 $Y=1177678
X85 401 16062 26 25 16174 NOR2BX1 $T=1541920 1325530 0 0 $X=1541918 $Y=1325278
X86 370 16185 26 25 16125 NOR2BX1 $T=1543760 1259110 1 180 $X=1541920 $Y=1258858
X87 401 16115 26 25 16119 NOR2BX1 $T=1544680 1303390 0 180 $X=1542840 $Y=1299450
X88 546 16185 26 25 16197 NOR2BX1 $T=1544220 1266490 1 0 $X=1544218 $Y=1262550
X89 536 16199 26 25 16124 NOR2BX1 $T=1546060 1192690 1 180 $X=1544220 $Y=1192438
X90 536 16188 26 25 16304 NOR2BX1 $T=1546980 1229590 0 0 $X=1546978 $Y=1229338
X91 546 16115 26 25 16221 NOR2BX1 $T=1549740 1303390 0 180 $X=1547900 $Y=1299450
X92 378 16246 26 25 16252 NOR2BX1 $T=1548820 1170550 1 0 $X=1548818 $Y=1166610
X93 364 16199 26 25 16231 NOR2BX1 $T=1550660 1192690 0 180 $X=1548820 $Y=1188750
X94 398 16213 26 25 16288 NOR2BX1 $T=1549740 1200070 0 0 $X=1549738 $Y=1199818
X95 546 16062 26 25 16273 NOR2BX1 $T=1549740 1325530 1 0 $X=1549738 $Y=1321590
X96 398 16293 26 25 16249 NOR2BX1 $T=1551580 1185310 1 180 $X=1549740 $Y=1185058
X97 536 16213 26 25 16171 NOR2BX1 $T=1551580 1214830 0 180 $X=1549740 $Y=1210890
X98 375 16092 26 25 16228 NOR2BX1 $T=1552500 1177930 1 180 $X=1550660 $Y=1177678
X99 364 16289 26 25 16298 NOR2BX1 $T=1552960 1310770 1 0 $X=1552958 $Y=1306830
X100 536 16246 26 25 16211 NOR2BX1 $T=1555720 1177930 0 180 $X=1553880 $Y=1173990
X101 546 16290 26 25 16299 NOR2BX1 $T=1555720 1347670 0 180 $X=1553880 $Y=1343730
X102 370 16356 26 25 16297 NOR2BX1 $T=1556180 1266490 1 180 $X=1554340 $Y=1266238
X103 536 16293 26 25 16326 NOR2BX1 $T=1555260 1185310 1 0 $X=1555258 $Y=1181370
X104 368 16290 26 25 16308 NOR2BX1 $T=1558020 1347670 0 180 $X=1556180 $Y=1343730
X105 458 16188 26 25 16307 NOR2BX1 $T=1560780 1229590 1 180 $X=1558940 $Y=1229338
X106 536 16359 26 25 16302 NOR2BX1 $T=1560780 1244350 1 180 $X=1558940 $Y=1244098
X107 546 16289 26 25 16395 NOR2BX1 $T=1560320 1310770 1 0 $X=1560318 $Y=1306830
X108 398 16386 26 25 16301 NOR2BX1 $T=1562160 1214830 1 180 $X=1560320 $Y=1214578
X109 485 16359 26 25 16319 NOR2BX1 $T=1562160 1251730 1 180 $X=1560320 $Y=1251478
X110 375 16393 26 25 16401 NOR2BX1 $T=1561700 1281250 0 0 $X=1561698 $Y=1280998
X111 398 16411 26 25 16348 NOR2BX1 $T=1564000 1185310 1 180 $X=1562160 $Y=1185058
X112 536 16356 26 25 16407 NOR2BX1 $T=1568140 1266490 1 180 $X=1566300 $Y=1266238
X113 536 16446 26 25 16467 NOR2BX1 $T=1567220 1177930 0 0 $X=1567218 $Y=1177678
X114 536 16386 26 25 16447 NOR2BX1 $T=1567220 1222210 1 0 $X=1567218 $Y=1218270
X115 536 16411 26 25 16416 NOR2BX1 $T=1573200 1192690 0 180 $X=1571360 $Y=1188750
X116 401 16446 26 25 16489 NOR2BX1 $T=1572740 1177930 0 0 $X=1572738 $Y=1177678
X117 546 16393 26 25 16487 NOR2BX1 $T=1574580 1288630 0 180 $X=1572740 $Y=1284690
X118 8881 25 8940 26 CLKBUFX3 $T=1060300 1192690 1 0 $X=1060298 $Y=1188750
X119 9006 25 8947 26 CLKBUFX3 $T=1070880 1192690 0 180 $X=1069040 $Y=1188750
X120 9225 25 8936 26 CLKBUFX3 $T=1085600 1185310 0 180 $X=1083760 $Y=1181370
X121 9380 25 32 26 CLKBUFX3 $T=1094800 1296010 0 0 $X=1094798 $Y=1295758
X122 50 25 9380 26 CLKBUFX3 $T=1104920 1303390 1 180 $X=1103080 $Y=1303138
X123 32 25 9644 26 CLKBUFX3 $T=1104460 1281250 1 0 $X=1104458 $Y=1277310
X124 9392 25 9532 26 CLKBUFX3 $T=1110440 1111510 0 0 $X=1110438 $Y=1111258
X125 32 25 9815 26 CLKBUFX3 $T=1114580 1251730 0 0 $X=1114578 $Y=1251478
X126 9791 25 9740 26 CLKBUFX3 $T=1115960 1170550 0 0 $X=1115958 $Y=1170298
X127 9851 25 9686 26 CLKBUFX3 $T=1119180 1296010 0 180 $X=1117340 $Y=1292070
X128 9363 25 9573 26 CLKBUFX3 $T=1121480 1104130 0 0 $X=1121478 $Y=1103878
X129 10231 25 8883 26 CLKBUFX3 $T=1136660 1259110 0 180 $X=1134820 $Y=1255170
X130 10297 25 8748 26 CLKBUFX3 $T=1139880 1251730 1 180 $X=1138040 $Y=1251478
X131 10310 25 8749 26 CLKBUFX3 $T=1140800 1229590 0 180 $X=1138960 $Y=1225650
X132 10312 25 10362 26 CLKBUFX3 $T=1139420 1288630 0 0 $X=1139418 $Y=1288378
X133 10364 25 8961 26 CLKBUFX3 $T=1142640 1222210 1 180 $X=1140800 $Y=1221958
X134 10382 25 9101 26 CLKBUFX3 $T=1144940 1185310 1 180 $X=1143100 $Y=1185058
X135 10291 25 10445 26 CLKBUFX3 $T=1144480 1288630 0 0 $X=1144478 $Y=1288378
X136 10409 25 8736 26 CLKBUFX3 $T=1144940 1251730 0 0 $X=1144938 $Y=1251478
X137 10413 25 8871 26 CLKBUFX3 $T=1145860 1259110 1 0 $X=1145858 $Y=1255170
X138 10292 25 10004 26 CLKBUFX3 $T=1149080 1288630 0 0 $X=1149078 $Y=1288378
X139 10556 25 9003 26 CLKBUFX3 $T=1152760 1185310 0 180 $X=1150920 $Y=1181370
X140 10260 25 10380 26 CLKBUFX3 $T=1151380 1266490 1 0 $X=1151378 $Y=1262550
X141 10640 25 8742 26 CLKBUFX3 $T=1156900 1251730 0 0 $X=1156898 $Y=1251478
X142 10617 25 8732 26 CLKBUFX3 $T=1156900 1266490 1 0 $X=1156898 $Y=1262550
X143 10657 25 85 26 CLKBUFX3 $T=1159200 1340290 1 180 $X=1157360 $Y=1340038
X144 9991 25 9729 26 CLKBUFX3 $T=1157820 1185310 1 0 $X=1157818 $Y=1181370
X145 10673 25 9102 26 CLKBUFX3 $T=1159660 1177930 1 180 $X=1157820 $Y=1177678
X146 125 25 10716 26 CLKBUFX3 $T=1158280 1288630 0 0 $X=1158278 $Y=1288378
X147 9729 25 9765 26 CLKBUFX3 $T=1161040 1155790 1 0 $X=1161038 $Y=1151850
X148 10470 25 10755 26 CLKBUFX3 $T=1161960 1074610 0 0 $X=1161958 $Y=1074358
X149 10751 25 10125 26 CLKBUFX3 $T=1163800 1266490 0 180 $X=1161960 $Y=1262550
X150 9624 25 9708 26 CLKBUFX3 $T=1162420 1148410 1 0 $X=1162418 $Y=1144470
X151 10528 25 10751 26 CLKBUFX3 $T=1162420 1273870 0 0 $X=1162418 $Y=1273618
X152 10605 25 10207 26 CLKBUFX3 $T=1163800 1126270 1 0 $X=1163798 $Y=1122330
X153 9920 25 10484 26 CLKBUFX3 $T=1163800 1148410 0 0 $X=1163798 $Y=1148158
X154 10758 25 8814 26 CLKBUFX3 $T=1164260 1236970 1 0 $X=1164258 $Y=1233030
X155 10813 25 8816 26 CLKBUFX3 $T=1166560 1244350 1 180 $X=1164720 $Y=1244098
X156 9196 25 10887 26 CLKBUFX3 $T=1167020 1126270 0 0 $X=1167018 $Y=1126018
X157 10469 25 10871 26 CLKBUFX3 $T=1168400 1148410 1 0 $X=1168398 $Y=1144470
X158 10893 25 9228 26 CLKBUFX3 $T=1170700 1222210 0 180 $X=1168860 $Y=1218270
X159 147 25 10184 26 CLKBUFX3 $T=1173920 1325530 1 180 $X=1172080 $Y=1325278
X160 10953 25 9270 26 CLKBUFX3 $T=1174380 1192690 1 180 $X=1172540 $Y=1192438
X161 10619 25 10951 26 CLKBUFX3 $T=1173000 1081990 1 0 $X=1172998 $Y=1078050
X162 10470 25 10750 26 CLKBUFX3 $T=1173920 1148410 1 0 $X=1173918 $Y=1144470
X163 9196 25 10908 26 CLKBUFX3 $T=1178060 1148410 1 0 $X=1178058 $Y=1144470
X164 10988 25 11052 26 CLKBUFX3 $T=1178060 1273870 1 0 $X=1178058 $Y=1269930
X165 147 25 138 26 CLKBUFX3 $T=1180820 1318150 1 180 $X=1178980 $Y=1317898
X166 9196 25 11133 26 CLKBUFX3 $T=1190480 1081990 1 0 $X=1190478 $Y=1078050
X167 147 25 99 26 CLKBUFX3 $T=1191860 1318150 0 0 $X=1191858 $Y=1317898
X168 11357 25 9386 26 CLKBUFX3 $T=1194160 1200070 0 180 $X=1192320 $Y=1196130
X169 10619 25 10299 26 CLKBUFX3 $T=1200140 1089370 0 180 $X=1198300 $Y=1085430
X170 10605 25 11030 26 CLKBUFX3 $T=1201980 1081990 0 0 $X=1201978 $Y=1081738
X171 11626 25 11706 26 CLKBUFX3 $T=1207960 1318150 0 0 $X=1207958 $Y=1317898
X172 11731 25 11736 26 CLKBUFX3 $T=1212560 1325530 1 0 $X=1212558 $Y=1321590
X173 10961 25 11899 26 CLKBUFX3 $T=1214400 1340290 1 0 $X=1214398 $Y=1336350
X174 201 25 11426 26 CLKBUFX3 $T=1216240 1296010 0 0 $X=1216238 $Y=1295758
X175 11992 25 12117 26 CLKBUFX3 $T=1227280 1325530 1 0 $X=1227278 $Y=1321590
X176 12155 25 11568 26 CLKBUFX3 $T=1233720 1281250 1 180 $X=1231880 $Y=1280998
X177 12172 25 11586 26 CLKBUFX3 $T=1234640 1332910 0 180 $X=1232800 $Y=1328970
X178 12172 25 12296 26 CLKBUFX3 $T=1241540 1332910 1 0 $X=1241538 $Y=1328970
X179 12352 25 12336 26 CLKBUFX3 $T=1243840 1325530 1 180 $X=1242000 $Y=1325278
X180 12358 25 12015 26 CLKBUFX3 $T=1244300 1259110 0 180 $X=1242460 $Y=1255170
X181 9840 25 9988 26 CLKBUFX3 $T=1243380 1067230 0 0 $X=1243378 $Y=1066978
X182 12144 25 12016 26 CLKBUFX3 $T=1244300 1273870 0 0 $X=1244298 $Y=1273618
X183 147 25 11850 26 CLKBUFX3 $T=1247520 1244350 0 0 $X=1247518 $Y=1244098
X184 12155 25 12270 26 CLKBUFX3 $T=1249820 1281250 0 0 $X=1249818 $Y=1280998
X185 50 25 281 26 CLKBUFX3 $T=1270980 1347670 1 0 $X=1270978 $Y=1343730
X186 281 25 201 26 CLKBUFX3 $T=1290760 1318150 0 180 $X=1288920 $Y=1314210
X187 13566 25 13646 26 CLKBUFX3 $T=1304560 1259110 1 0 $X=1304558 $Y=1255170
X188 13726 25 67 26 CLKBUFX3 $T=1313760 1347670 0 180 $X=1311920 $Y=1343730
X189 39 25 13981 26 CLKBUFX3 $T=1333080 1340290 0 0 $X=1333078 $Y=1340038
X190 13981 25 13883 26 CLKBUFX3 $T=1349180 1310770 1 0 $X=1349178 $Y=1306830
X191 14150 25 348 26 CLKBUFX3 $T=1351940 1340290 1 0 $X=1351938 $Y=1336350
X192 53 25 430 26 CLKBUFX3 $T=1367580 1192690 1 0 $X=1367578 $Y=1188750
X193 83 25 425 26 CLKBUFX3 $T=1374480 1214830 0 0 $X=1374478 $Y=1214578
X194 454 25 14191 26 CLKBUFX3 $T=1390580 1244350 1 0 $X=1390578 $Y=1240410
X195 452 25 14639 26 CLKBUFX3 $T=1398860 1340290 0 0 $X=1398858 $Y=1340038
X196 281 25 466 26 CLKBUFX3 $T=1404840 1347670 0 0 $X=1404838 $Y=1347418
X197 14732 25 14837 26 CLKBUFX3 $T=1410360 1214830 1 0 $X=1410358 $Y=1210890
X198 450 25 474 26 CLKBUFX3 $T=1414960 1347670 1 0 $X=1414958 $Y=1343730
X199 281 25 362 26 CLKBUFX3 $T=1416340 1340290 0 0 $X=1416338 $Y=1340038
X200 12142 25 14913 26 CLKBUFX3 $T=1420020 1126270 1 0 $X=1420018 $Y=1122330
X201 12063 25 14867 26 CLKBUFX3 $T=1420940 1111510 0 0 $X=1420938 $Y=1111258
X202 12024 25 14926 26 CLKBUFX3 $T=1420940 1310770 0 0 $X=1420938 $Y=1310518
X203 479 25 352 26 CLKBUFX3 $T=1420940 1332910 0 0 $X=1420938 $Y=1332658
X204 12039 25 14879 26 CLKBUFX3 $T=1421860 1222210 1 0 $X=1421858 $Y=1218270
X205 454 25 422 26 CLKBUFX3 $T=1421860 1325530 1 0 $X=1421858 $Y=1321590
X206 12050 25 14917 26 CLKBUFX3 $T=1423700 1266490 1 0 $X=1423698 $Y=1262550
X207 12051 25 14937 26 CLKBUFX3 $T=1428760 1288630 0 0 $X=1428758 $Y=1288378
X208 12792 25 14993 26 CLKBUFX3 $T=1429220 1111510 1 0 $X=1429218 $Y=1107570
X209 12143 25 14955 26 CLKBUFX3 $T=1431980 1192690 0 0 $X=1431978 $Y=1192438
X210 490 25 13915 26 CLKBUFX3 $T=1432440 1266490 1 0 $X=1432438 $Y=1262550
X211 490 25 495 26 CLKBUFX3 $T=1432440 1266490 0 0 $X=1432438 $Y=1266238
X212 12110 25 15022 26 CLKBUFX3 $T=1432440 1318150 1 0 $X=1432438 $Y=1314210
X213 78 25 410 26 CLKBUFX3 $T=1432900 1236970 0 0 $X=1432898 $Y=1236718
X214 479 25 13880 26 CLKBUFX3 $T=1433360 1229590 0 0 $X=1433358 $Y=1229338
X215 13390 25 15053 26 CLKBUFX3 $T=1437500 1259110 0 0 $X=1437498 $Y=1258858
X216 479 25 361 26 CLKBUFX3 $T=1438420 1318150 1 0 $X=1438418 $Y=1314210
X217 78 25 426 26 CLKBUFX3 $T=1438880 1251730 1 0 $X=1438878 $Y=1247790
X218 12516 25 15020 26 CLKBUFX3 $T=1439340 1118890 1 0 $X=1439338 $Y=1114950
X219 12258 25 14929 26 CLKBUFX3 $T=1439340 1332910 1 0 $X=1439338 $Y=1328970
X220 493 25 15075 26 CLKBUFX3 $T=1440720 1296010 1 0 $X=1440718 $Y=1292070
X221 489 25 14921 26 CLKBUFX3 $T=1442100 1273870 0 0 $X=1442098 $Y=1273618
X222 495 25 354 26 CLKBUFX3 $T=1442560 1273870 1 0 $X=1442558 $Y=1269930
X223 495 25 14119 26 CLKBUFX3 $T=1443480 1207450 1 0 $X=1443478 $Y=1203510
X224 12754 25 14992 26 CLKBUFX3 $T=1444400 1118890 1 0 $X=1444398 $Y=1114950
X225 424 25 429 26 CLKBUFX3 $T=1446240 1266490 0 0 $X=1446238 $Y=1266238
X226 496 25 14936 26 CLKBUFX3 $T=1447160 1273870 1 0 $X=1447158 $Y=1269930
X227 12589 25 14966 26 CLKBUFX3 $T=1449460 1111510 1 0 $X=1449458 $Y=1107570
X228 13329 25 15224 26 CLKBUFX3 $T=1451300 1273870 1 0 $X=1451298 $Y=1269930
X229 385 25 387 26 CLKBUFX3 $T=1451760 1236970 0 0 $X=1451758 $Y=1236718
X230 495 25 13853 26 CLKBUFX3 $T=1460960 1325530 0 0 $X=1460958 $Y=1325278
X231 495 25 366 26 CLKBUFX3 $T=1462800 1296010 1 0 $X=1462798 $Y=1292070
X232 518 25 513 26 CLKBUFX3 $T=1466940 1325530 0 180 $X=1465100 $Y=1321590
X233 521 25 381 26 CLKBUFX3 $T=1470160 1259110 0 180 $X=1468320 $Y=1255170
X234 495 25 13893 26 CLKBUFX3 $T=1468780 1318150 1 0 $X=1468778 $Y=1314210
X235 13883 25 14264 26 CLKBUFX3 $T=1469240 1244350 1 0 $X=1469238 $Y=1240410
X236 13405 25 15427 26 CLKBUFX3 $T=1473380 1229590 0 0 $X=1473378 $Y=1229338
X237 514 25 15057 26 CLKBUFX3 $T=1475680 1281250 1 0 $X=1475678 $Y=1277310
X238 521 25 14098 26 CLKBUFX3 $T=1477980 1207450 1 180 $X=1476140 $Y=1207198
X239 521 25 371 26 CLKBUFX3 $T=1477520 1229590 0 0 $X=1477518 $Y=1229338
X240 13332 25 15523 26 CLKBUFX3 $T=1481660 1229590 0 0 $X=1481658 $Y=1229338
X241 78 25 413 26 CLKBUFX3 $T=1485800 1229590 0 0 $X=1485798 $Y=1229338
X242 506 25 15131 26 CLKBUFX3 $T=1486260 1288630 1 0 $X=1486258 $Y=1284690
X243 15292 25 15437 26 CLKBUFX3 $T=1486260 1296010 1 0 $X=1486258 $Y=1292070
X244 517 25 15296 26 CLKBUFX3 $T=1487180 1281250 1 0 $X=1487178 $Y=1277310
X245 520 25 15253 26 CLKBUFX3 $T=1489480 1288630 1 0 $X=1489478 $Y=1284690
X246 535 25 369 26 CLKBUFX3 $T=1494080 1266490 1 0 $X=1494078 $Y=1262550
X247 526 25 15352 26 CLKBUFX3 $T=1506500 1296010 0 180 $X=1504660 $Y=1292070
X248 521 25 13891 26 CLKBUFX3 $T=1509260 1185310 0 180 $X=1507420 $Y=1181370
X249 546 25 530 26 CLKBUFX3 $T=1508340 1347670 1 0 $X=1508338 $Y=1343730
X250 14732 25 15353 26 CLKBUFX3 $T=1509260 1200070 0 0 $X=1509258 $Y=1199818
X251 495 25 13879 26 CLKBUFX3 $T=1511560 1192690 1 180 $X=1509720 $Y=1192438
X252 521 25 13912 26 CLKBUFX3 $T=1511560 1332910 1 180 $X=1509720 $Y=1332658
X253 14264 25 551 26 CLKBUFX3 $T=1514780 1281250 0 0 $X=1514778 $Y=1280998
X254 533 25 15313 26 CLKBUFX3 $T=1514780 1296010 0 0 $X=1514778 $Y=1295758
X255 15631 25 15760 26 CLKBUFX3 $T=1517080 1318150 1 180 $X=1515240 $Y=1317898
X256 529 25 15439 26 CLKBUFX3 $T=1519840 1296010 0 0 $X=1519838 $Y=1295758
X257 90 25 536 26 CLKBUFX3 $T=1520760 1347670 0 0 $X=1520758 $Y=1347418
X258 550 25 412 26 CLKBUFX3 $T=1523060 1325530 0 0 $X=1523058 $Y=1325278
X259 495 25 360 26 CLKBUFX3 $T=1525360 1340290 1 180 $X=1523520 $Y=1340038
X260 318 25 548 26 CLKBUFX3 $T=1523980 1347670 0 0 $X=1523978 $Y=1347418
X261 550 25 535 26 CLKBUFX3 $T=1524900 1340290 1 0 $X=1524898 $Y=1336350
X262 550 25 373 26 CLKBUFX3 $T=1525820 1332910 0 0 $X=1525818 $Y=1332658
X263 281 25 15996 26 CLKBUFX3 $T=1527200 1347670 0 0 $X=1527198 $Y=1347418
X264 495 25 365 26 CLKBUFX3 $T=1529040 1347670 0 180 $X=1527200 $Y=1343730
X265 550 25 415 26 CLKBUFX3 $T=1527660 1340290 0 0 $X=1527658 $Y=1340038
X266 495 25 561 26 CLKBUFX3 $T=1530420 1251730 1 0 $X=1530418 $Y=1247790
X267 562 25 15631 26 CLKBUFX3 $T=1532260 1325530 1 0 $X=1532258 $Y=1321590
X268 550 25 13974 26 CLKBUFX3 $T=1536860 1325530 0 0 $X=1536858 $Y=1325278
X269 550 25 389 26 CLKBUFX3 $T=1537320 1332910 1 0 $X=1537318 $Y=1328970
X270 557 25 568 26 CLKBUFX3 $T=1537320 1347670 0 0 $X=1537318 $Y=1347418
X271 521 25 16095 26 CLKBUFX3 $T=1544220 1318150 0 0 $X=1544218 $Y=1317898
X272 495 25 567 26 CLKBUFX3 $T=1544680 1281250 0 0 $X=1544678 $Y=1280998
X273 587 25 586 26 CLKBUFX3 $T=1563540 1318150 1 180 $X=1561700 $Y=1317898
X274 562 25 15942 26 CLKBUFX3 $T=1587920 1288630 0 0 $X=1587918 $Y=1288378
X275 16449 25 76 26 CLKBUFX3 $T=1587920 1318150 0 0 $X=1587918 $Y=1317898
X276 16720 25 9816 26 CLKBUFX3 $T=1598960 1318150 1 180 $X=1597120 $Y=1317898
X277 16720 25 16449 26 CLKBUFX3 $T=1601720 1318150 1 0 $X=1601718 $Y=1314210
X278 50 25 16720 26 CLKBUFX3 $T=1607240 1318150 1 0 $X=1607238 $Y=1314210
X279 16720 25 622 26 CLKBUFX3 $T=1608160 1325530 1 0 $X=1608158 $Y=1321590
X280 9519 9382 9382 25 9430 26 9622 OAI2BB2XL $T=1102620 1310770 0 0 $X=1102618 $Y=1310518
X281 51 16400 16414 25 16421 26 16434 OAI2BB2XL $T=1562620 1273870 0 0 $X=1562618 $Y=1273618
X282 87 16442 16400 25 16444 26 16515 OAI2BB2XL $T=1565380 1244350 0 0 $X=1565378 $Y=1244098
X283 264 16485 599 25 16482 26 16428 OAI2BB2XL $T=1573660 1340290 0 180 $X=1570900 $Y=1336350
X284 55 16442 16414 25 16413 26 16518 OAI2BB2XL $T=1571360 1251730 0 0 $X=1571358 $Y=1251478
X285 143 16442 16414 25 16495 26 16453 OAI2BB2XL $T=1571820 1214830 0 0 $X=1571818 $Y=1214578
X286 40 16400 16400 25 16496 26 16427 OAI2BB2XL $T=1571820 1310770 1 0 $X=1571818 $Y=1306830
X287 289 16442 16414 25 16438 26 16514 OAI2BB2XL $T=1572740 1236970 1 0 $X=1572738 $Y=1233030
X288 100 16400 16400 25 16510 26 16525 OAI2BB2XL $T=1572740 1244350 1 0 $X=1572738 $Y=1240410
X289 227 16400 604 25 598 26 16529 OAI2BB2XL $T=1579180 1318150 1 180 $X=1576420 $Y=1317898
X290 70 16400 16414 25 16543 26 16547 OAI2BB2XL $T=1576880 1296010 1 0 $X=1576878 $Y=1292070
X291 308 16442 16414 25 16545 26 16563 OAI2BB2XL $T=1577340 1266490 1 0 $X=1577338 $Y=1262550
X292 56 16400 16400 25 16546 26 16564 OAI2BB2XL $T=1577340 1273870 1 0 $X=1577338 $Y=1269930
X293 45 16400 16485 25 16552 26 16540 OAI2BB2XL $T=1577800 1303390 1 0 $X=1577798 $Y=1299450
X294 109 16400 16400 25 16541 26 16598 OAI2BB2XL $T=1578720 1318150 1 0 $X=1578718 $Y=1314210
X295 124 16442 16414 25 16466 26 16612 OAI2BB2XL $T=1579180 1222210 1 0 $X=1579178 $Y=1218270
X296 111 16442 16400 25 16542 26 16538 OAI2BB2XL $T=1579180 1236970 0 0 $X=1579178 $Y=1236718
X297 241 16485 16400 25 16439 26 16548 OAI2BB2XL $T=1581940 1340290 0 180 $X=1579180 $Y=1336350
X298 177 16485 604 25 16568 26 16593 OAI2BB2XL $T=1579640 1318150 0 0 $X=1579638 $Y=1317898
X299 80 16400 16414 25 16581 26 16539 OAI2BB2XL $T=1580100 1251730 0 0 $X=1580098 $Y=1251478
X300 139 16442 16414 25 16626 26 16771 OAI2BB2XL $T=1587920 1222210 1 0 $X=1587918 $Y=1218270
X301 300 16442 16414 25 16627 26 16582 OAI2BB2XL $T=1587920 1273870 0 0 $X=1587918 $Y=1273618
X302 75 16400 16414 25 16362 26 16605 OAI2BB2XL $T=1592520 1259110 1 180 $X=1589760 $Y=1258858
X303 213 16400 604 25 16602 26 16588 OAI2BB2XL $T=1592520 1310770 0 180 $X=1589760 $Y=1306830
X304 235 16485 604 25 16594 26 16632 OAI2BB2XL $T=1592520 1325530 1 180 $X=1589760 $Y=1325278
X305 280 16442 16414 25 16645 26 16723 OAI2BB2XL $T=1594360 1288630 0 0 $X=1594358 $Y=1288378
X306 231 16485 604 25 16646 26 16697 OAI2BB2XL $T=1594360 1332910 1 0 $X=1594358 $Y=1328970
X307 616 16442 16414 25 16692 26 16691 OAI2BB2XL $T=1597120 1259110 1 180 $X=1594360 $Y=1258858
X308 618 16442 16442 25 16693 26 16673 OAI2BB2XL $T=1597120 1273870 0 180 $X=1594360 $Y=1269930
X309 309 16485 604 25 16719 26 16674 OAI2BB2XL $T=1596200 1296010 0 0 $X=1596198 $Y=1295758
X310 621 619 604 25 16620 26 16589 OAI2BB2XL $T=1599420 1347670 1 180 $X=1596660 $Y=1347418
X311 284 16485 604 25 16684 26 16711 OAI2BB2XL $T=1599880 1310770 0 180 $X=1597120 $Y=1306830
X312 242 16485 604 25 16703 26 16733 OAI2BB2XL $T=1603560 1325530 1 180 $X=1600800 $Y=1325278
X313 321 16442 16414 25 16600 26 16731 OAI2BB2XL $T=1604480 1266490 1 180 $X=1601720 $Y=1266238
X314 279 16442 16414 25 16714 26 16775 OAI2BB2XL $T=1604020 1229590 0 0 $X=1604018 $Y=1229338
X315 623 16442 16414 25 16702 26 16769 OAI2BB2XL $T=1607240 1266490 0 180 $X=1604480 $Y=1262550
X316 624 16400 16414 25 16683 26 16770 OAI2BB2XL $T=1607240 1288630 0 180 $X=1604480 $Y=1284690
X317 628 16485 16485 25 16688 26 16766 OAI2BB2XL $T=1608160 1296010 1 180 $X=1605400 $Y=1295758
X318 629 619 604 25 16554 26 16624 OAI2BB2XL $T=1608160 1347670 1 180 $X=1605400 $Y=1347418
X319 117 16442 16400 25 16765 26 16690 OAI2BB2XL $T=1609540 1244350 1 180 $X=1606780 $Y=1244098
X320 631 16825 604 25 16768 26 16821 OAI2BB2XL $T=1614140 1310770 0 180 $X=1611380 $Y=1306830
X321 639 16485 16414 25 16783 26 16732 OAI2BB2XL $T=1615980 1288630 1 180 $X=1613220 $Y=1288378
X322 632 16442 16414 25 16778 26 16830 OAI2BB2XL $T=1617360 1273870 0 180 $X=1614600 $Y=1269930
X323 635 16825 16825 25 16831 26 16829 OAI2BB2XL $T=1617360 1332910 1 180 $X=1614600 $Y=1332658
X324 634 16825 16825 25 16763 26 16819 OAI2BB2XL $T=1621500 1296010 1 180 $X=1618740 $Y=1295758
X325 643 16825 604 25 16832 26 16880 OAI2BB2XL $T=1624720 1340290 0 180 $X=1621960 $Y=1336350
X326 637 16442 16414 25 16767 26 16822 OAI2BB2XL $T=1626100 1281250 0 180 $X=1623340 $Y=1277310
X327 641 16825 604 25 16823 26 16847 OAI2BB2XL $T=1627020 1325530 1 180 $X=1624260 $Y=1325278
X328 642 625 604 25 16824 26 16848 OAI2BB2XL $T=1627020 1347670 0 180 $X=1624260 $Y=1343730
X329 640 16825 16825 25 16820 26 16879 OAI2BB2XL $T=1627480 1303390 1 180 $X=1624720 $Y=1303138
X330 644 16825 16825 25 16834 26 16886 OAI2BB2XL $T=1627480 1318150 0 180 $X=1624720 $Y=1314210
X331 638 16825 16825 25 16762 26 16826 OAI2BB2XL $T=1627940 1310770 1 180 $X=1625180 $Y=1310518
X332 550 376 25 26 CLKBUFX4 $T=1525360 1340290 0 0 $X=1525358 $Y=1340038
X333 550 386 25 26 CLKBUFX4 $T=1542380 1332910 1 0 $X=1542378 $Y=1328970
X334 9069 29 9072 30 32 33 26 25 36 SDFFRXL $T=1074100 1347670 0 0 $X=1074098 $Y=1347418
X335 9069 9213 9202 30 32 9072 26 25 28 SDFFRXL $T=1085140 1340290 0 180 $X=1074100 $Y=1336350
X336 9069 9523 9511 9404 32 9351 26 25 9336 SDFFRXL $T=1104000 1259110 1 180 $X=1092960 $Y=1258858
X337 9069 9524 9336 9404 32 9340 26 25 9337 SDFFRXL $T=1104000 1281250 0 180 $X=1092960 $Y=1277310
X338 9069 9361 9378 9404 32 9541 26 25 9511 SDFFRXL $T=1093420 1266490 1 0 $X=1093418 $Y=1262550
X339 9069 9372 40 9404 32 9554 26 25 9576 SDFFRXL $T=1093880 1281250 0 0 $X=1093878 $Y=1280998
X340 9069 9594 9337 9404 9557 9418 26 25 9398 SDFFRXL $T=1107220 1273870 1 180 $X=1096180 $Y=1273618
X341 9069 9616 51 9404 32 9371 26 25 9408 SDFFRXL $T=1107680 1259110 0 180 $X=1096640 $Y=1255170
X342 9069 9617 56 9404 32 9425 26 25 9378 SDFFRXL $T=1107680 1266490 1 180 $X=1096640 $Y=1266238
X343 9069 9622 9595 9404 32 9430 26 25 9421 SDFFRXL $T=1108140 1310770 0 180 $X=1097100 $Y=1306830
X344 9069 9623 9421 30 32 9431 26 25 9405 SDFFRXL $T=1108140 1318150 0 180 $X=1097100 $Y=1314210
X345 9069 9365 9431 30 50 9274 26 25 9419 SDFFRXL $T=1097560 1325530 1 0 $X=1097558 $Y=1321590
X346 9069 9744 9722 9404 32 9553 26 25 9526 SDFFRXL $T=1114580 1251730 1 180 $X=1103540 $Y=1251478
X347 9664 61 62 30 76 9861 26 25 82 SDFFRXL $T=1108600 1347670 0 0 $X=1108598 $Y=1347418
X348 9069 9848 9828 9404 9557 9395 26 25 9655 SDFFRXL $T=1119640 1273870 1 180 $X=1108600 $Y=1273618
X349 9664 9682 9706 30 9816 9804 26 25 9931 SDFFRXL $T=1109520 1332910 1 0 $X=1109518 $Y=1328970
X350 9069 9738 9655 9404 9557 9903 26 25 95 SDFFRXL $T=1111820 1288630 1 0 $X=1111818 $Y=1284690
X351 9664 9669 9792 30 9816 9706 26 25 10104 SDFFRXL $T=1113660 1340290 1 0 $X=1113658 $Y=1336350
X352 9780 9781 9786 9404 9815 9974 26 25 9996 SDFFRXL $T=1114120 1229590 0 0 $X=1114118 $Y=1229338
X353 9664 9783 9804 30 9816 9976 26 25 9705 SDFFRXL $T=1114120 1325530 1 0 $X=1114118 $Y=1321590
X354 9069 9966 9408 9404 9815 9699 26 25 9767 SDFFRXL $T=1125160 1259110 1 180 $X=1114120 $Y=1258858
X355 9069 9967 45 9404 9644 9782 26 25 9768 SDFFRXL $T=1125160 1281250 0 180 $X=1114120 $Y=1277310
X356 9780 9975 87 9404 9815 9721 26 25 9722 SDFFRXL $T=1125620 1244350 0 180 $X=1114580 $Y=1240410
X357 9664 9977 9861 30 76 9792 26 25 9776 SDFFRXL $T=1125620 1340290 1 180 $X=1114580 $Y=1340038
X358 9780 9801 75 9404 9815 10003 26 25 10020 SDFFRXL $T=1115040 1229590 1 0 $X=1115038 $Y=1225650
X359 9780 9992 9964 9404 9815 9802 26 25 9662 SDFFRXL $T=1126080 1244350 1 180 $X=1115040 $Y=1244098
X360 9780 9993 55 9404 9815 9763 26 25 9786 SDFFRXL $T=1126080 1251730 0 180 $X=1115040 $Y=1247790
X361 9780 10031 80 9404 9815 10238 26 25 10219 SDFFRXL $T=1126080 1214830 0 0 $X=1126078 $Y=1214578
X362 9780 10237 10219 9404 9815 10039 26 25 10025 SDFFRXL $T=1137580 1214830 0 180 $X=1126540 $Y=1210890
X363 9664 10249 10103 30 10184 10041 26 25 10033 SDFFRXL $T=1138040 1332910 0 180 $X=1127000 $Y=1328970
X364 9664 10256 10041 30 10184 10054 26 25 10035 SDFFRXL $T=1138500 1325530 1 180 $X=1127460 $Y=1325278
X365 9664 10293 10271 30 99 10103 26 25 10082 SDFFRXL $T=1140340 1332910 1 180 $X=1129300 $Y=1332658
X366 9664 10149 10157 30 10184 10301 26 25 10311 SDFFRXL $T=1130680 1318150 0 0 $X=1130678 $Y=1317898
X367 9664 10320 10301 9404 99 9595 26 25 10126 SDFFRXL $T=1141720 1310770 0 180 $X=1130680 $Y=1306830
X368 9780 10156 10152 9404 9815 10350 26 25 9964 SDFFRXL $T=1131140 1244350 0 0 $X=1131138 $Y=1244098
X369 9664 10335 10054 30 10184 10157 26 25 10044 SDFFRXL $T=1142180 1325530 0 180 $X=1131140 $Y=1321590
X370 9780 10351 109 9404 9815 10075 26 25 10152 SDFFRXL $T=1142640 1251730 0 180 $X=1131600 $Y=1247790
X371 9780 10361 10025 9404 9644 10063 26 25 10158 SDFFRXL $T=1143100 1200070 1 180 $X=1132060 $Y=1199818
X372 9780 10107 10198 9404 9815 10300 26 25 10390 SDFFRXL $T=1132520 1222210 1 0 $X=1132518 $Y=1218270
X373 9664 10543 9976 9404 50 10372 26 25 9470 SDFFRXL $T=1152300 1310770 1 180 $X=1141260 $Y=1310518
X374 9664 10488 10446 30 10184 10271 26 25 10354 SDFFRXL $T=1152300 1325530 1 180 $X=1141260 $Y=1325278
X375 9780 10401 111 9404 9644 10580 26 25 10198 SDFFRXL $T=1143100 1200070 1 0 $X=1143098 $Y=1196130
X376 10521 10269 117 9404 9815 10420 26 25 10229 SDFFRXL $T=1155520 1236970 0 180 $X=1144480 $Y=1233030
X377 10599 10440 10515 9404 10184 10422 26 25 10415 SDFFRXL $T=1155520 1303390 0 180 $X=1144480 $Y=1299450
X378 9664 120 10582 30 10184 10446 26 25 10430 SDFFRXL $T=1156440 1332910 0 180 $X=1145400 $Y=1328970
X379 9664 10437 10422 30 10184 10424 26 25 10487 SDFFRXL $T=1159200 1318150 0 180 $X=1148160 $Y=1314210
X380 10521 10352 70 9404 9815 10534 26 25 10683 SDFFRXL $T=1148620 1273870 1 0 $X=1148618 $Y=1269930
X381 9664 10522 10424 30 10184 10655 26 25 10705 SDFFRXL $T=1148620 1318150 0 0 $X=1148618 $Y=1317898
X382 9780 10448 124 9404 9644 10408 26 25 10439 SDFFRXL $T=1159660 1192690 1 180 $X=1148620 $Y=1192438
X383 9780 10532 10549 9404 9644 10703 26 25 10713 SDFFRXL $T=1149540 1185310 0 0 $X=1149538 $Y=1185058
X384 9780 10533 10158 9404 9644 10704 26 25 10714 SDFFRXL $T=1149540 1207450 0 0 $X=1149538 $Y=1207198
X385 10521 10449 100 9404 9815 10539 26 25 10645 SDFFRXL $T=1149540 1229590 0 0 $X=1149538 $Y=1229338
X386 9664 10736 10722 9404 10184 10581 26 25 10567 SDFFRXL $T=1163340 1310770 1 180 $X=1152300 $Y=1310518
X387 9664 10737 10655 30 10184 10582 26 25 10568 SDFFRXL $T=1163340 1325530 1 180 $X=1152300 $Y=1325278
X388 10599 10589 10581 9404 10184 10515 26 25 10596 SDFFRXL $T=1165180 1303390 1 180 $X=1154140 $Y=1303138
X389 10521 10905 10833 10868 9815 10734 26 25 10723 SDFFRXL $T=1172080 1251730 1 180 $X=1161040 $Y=1251478
X390 10521 10941 10780 10868 9557 10715 26 25 10757 SDFFRXL $T=1174380 1236970 1 180 $X=1163340 $Y=1236718
X391 10521 10950 10859 10868 9644 10768 26 25 9828 SDFFRXL $T=1174840 1273870 0 180 $X=1163800 $Y=1269930
X392 10521 10959 10940 9404 9815 10789 26 25 10780 SDFFRXL $T=1175300 1229590 0 180 $X=1164260 $Y=1225650
X393 9780 10981 139 9404 9557 10829 26 25 10812 SDFFRXL $T=1176680 1214830 0 180 $X=1165640 $Y=1210890
X394 10599 10841 10372 10868 9644 10960 26 25 11042 SDFFRXL $T=1166100 1303390 1 0 $X=1166098 $Y=1299450
X395 10599 10842 10858 10868 138 10795 26 25 10985 SDFFRXL $T=1166100 1310770 0 0 $X=1166098 $Y=1310518
X396 9780 10996 143 9404 9644 10765 26 25 10549 SDFFRXL $T=1177140 1192690 0 180 $X=1166100 $Y=1188750
X397 9780 10997 10812 9404 9644 10767 26 25 10823 SDFFRXL $T=1177140 1207450 0 180 $X=1166100 $Y=1203510
X398 10599 10801 10795 10868 138 10722 26 25 10824 SDFFRXL $T=1177140 1318150 0 180 $X=1166100 $Y=1314210
X399 10521 11006 10757 10868 9557 10808 26 25 10833 SDFFRXL $T=1177600 1244350 1 180 $X=1166560 $Y=1244098
X400 10521 11041 10723 10868 9557 10790 26 25 10859 SDFFRXL $T=1178980 1259110 1 180 $X=1167940 $Y=1258858
X401 10521 11022 11040 9404 9557 11129 26 25 10940 SDFFRXL $T=1175760 1229590 1 0 $X=1175758 $Y=1225650
X402 10599 11024 11042 10868 9644 11104 26 25 167 SDFFRXL $T=1175760 1303390 0 0 $X=1175758 $Y=1303138
X403 10521 11239 11221 9404 9815 11059 26 25 11040 SDFFRXL $T=1189100 1222210 1 180 $X=1178060 $Y=1221958
X404 9780 10837 174 9404 9644 11091 26 25 11084 SDFFRXL $T=1192320 1192690 0 180 $X=1181280 $Y=1188750
X405 10599 11304 11283 10868 11270 11137 26 25 10674 SDFFRXL $T=1192320 1310770 0 180 $X=1181280 $Y=1306830
X406 10599 11333 11137 10868 11270 10858 26 25 10612 SDFFRXL $T=1193700 1310770 1 180 $X=1182660 $Y=1310518
X407 9780 11154 10823 9404 9557 11352 26 25 11221 SDFFRXL $T=1183120 1207450 0 0 $X=1183118 $Y=1207198
X408 10599 11175 11195 10868 9557 11355 26 25 11364 SDFFRXL $T=1183120 1273870 0 0 $X=1183118 $Y=1273618
X409 10599 11267 11319 10868 11270 11174 26 25 10843 SDFFRXL $T=1194160 1266490 1 180 $X=1183120 $Y=1266238
X410 10599 11252 177 10868 9644 11123 26 25 11165 SDFFRXL $T=1194620 1296010 0 180 $X=1183580 $Y=1292070
X411 10599 11240 11165 10868 9644 11356 26 25 180 SDFFRXL $T=1186800 1303390 0 0 $X=1186798 $Y=1303138
X412 10599 11311 11174 10868 11270 11466 26 25 11282 SDFFRXL $T=1190480 1273870 1 0 $X=1190478 $Y=1269930
X413 11396 11402 11417 10868 11270 11418 26 25 10781 SDFFRXL $T=1195540 1244350 0 0 $X=1195538 $Y=1244098
X414 11396 179 11418 10868 11426 11319 26 25 10925 SDFFRXL $T=1195540 1259110 0 0 $X=1195538 $Y=1258858
X415 10521 188 11547 9404 11426 11395 26 25 10492 SDFFRXL $T=1206580 1207450 1 180 $X=1195540 $Y=1207198
X416 10599 189 11466 10868 11426 11409 26 25 11009 SDFFRXL $T=1207040 1266490 0 180 $X=1196000 $Y=1262550
X417 10599 11575 11491 10868 11270 11403 26 25 10849 SDFFRXL $T=1207040 1281250 1 180 $X=1196000 $Y=1280998
X418 11396 11562 11408 10868 11426 11407 26 25 11008 SDFFRXL $T=1207500 1236970 1 180 $X=1196460 $Y=1236718
X419 11396 11579 11409 10868 11270 11408 26 25 10973 SDFFRXL $T=1207500 1251730 1 180 $X=1196460 $Y=1251478
X420 11396 11246 11490 10868 11426 11417 26 25 10894 SDFFRXL $T=1208880 1244350 0 180 $X=1197840 $Y=1240410
X421 10599 11492 11403 10868 11270 11283 26 25 10769 SDFFRXL $T=1208880 1296010 1 180 $X=1197840 $Y=1295758
X422 10521 11315 11503 9404 11426 11547 26 25 11671 SDFFRXL $T=1199680 1200070 0 0 $X=1199678 $Y=1199818
X423 10521 195 11632 9404 11426 11490 26 25 10648 SDFFRXL $T=1211180 1229590 0 180 $X=1200140 $Y=1225650
X424 10599 196 11634 10868 11426 11491 26 25 10956 SDFFRXL $T=1211180 1296010 0 180 $X=1200140 $Y=1292070
X425 10521 11504 11395 9404 11426 11632 26 25 11430 SDFFRXL $T=1200600 1222210 0 0 $X=1200598 $Y=1221958
X426 10521 197 11644 9404 11426 11503 26 25 11442 SDFFRXL $T=1211640 1200070 0 180 $X=1200600 $Y=1196130
X427 11396 11522 11407 10868 11270 11704 26 25 10800 SDFFRXL $T=1201520 1236970 1 0 $X=1201518 $Y=1233030
X428 10521 11819 11870 11826 11850 11644 26 25 11415 SDFFRXL $T=1220380 1192690 1 180 $X=1209340 $Y=1192438
X429 11737 199 11753 10868 201 11939 26 25 10600 SDFFRXL $T=1212560 1332910 1 0 $X=1212558 $Y=1328970
X430 11737 210 11946 10868 201 11753 26 25 10558 SDFFRXL $T=1224980 1332910 1 180 $X=1213940 $Y=1332658
X431 11737 11993 11939 10868 99 11815 26 25 11086 SDFFRXL $T=1226360 1325530 0 180 $X=1215320 $Y=1321590
X432 11737 11868 213 10868 9644 11780 26 25 11195 SDFFRXL $T=1227740 1273870 1 180 $X=1216700 $Y=1273618
X433 11737 204 11815 10868 201 12052 26 25 10557 SDFFRXL $T=1217160 1310770 0 0 $X=1217158 $Y=1310518
X434 10521 216 11878 11826 11426 11870 26 25 11441 SDFFRXL $T=1228660 1192690 0 180 $X=1217620 $Y=1188750
X435 11737 217 12023 10868 11426 11634 26 25 10456 SDFFRXL $T=1228660 1296010 0 180 $X=1217620 $Y=1292070
X436 11737 203 11898 10868 201 12023 26 25 10641 SDFFRXL $T=1218080 1296010 0 0 $X=1218078 $Y=1295758
X437 10521 12062 12037 11826 11850 11878 26 25 11840 SDFFRXL $T=1229120 1200070 0 180 $X=1218080 $Y=1196130
X438 11737 12256 12052 10868 99 11898 26 25 11043 SDFFRXL $T=1240620 1303390 1 180 $X=1229580 $Y=1303138
X439 11396 12114 11704 11826 11270 12295 26 25 10730 SDFFRXL $T=1230040 1236970 1 0 $X=1230038 $Y=1233030
X440 11737 12297 12150 10868 99 11946 26 25 11604 SDFFRXL $T=1241540 1340290 1 180 $X=1230500 $Y=1340038
X441 12313 12303 12237 11826 11850 12037 26 25 12118 SDFFRXL $T=1242000 1200070 0 180 $X=1230960 $Y=1196130
X442 11737 12173 12213 10868 99 12150 26 25 11312 SDFFRXL $T=1242920 1347670 0 180 $X=1231880 $Y=1343730
X443 11396 12344 12295 10868 11850 12170 26 25 11410 SDFFRXL $T=1243840 1236970 1 180 $X=1232800 $Y=1236718
X444 233 232 12349 10868 99 12213 26 25 159 SDFFRXL $T=1245220 1347670 1 180 $X=1234180 $Y=1347418
X445 11396 12232 12216 10868 9644 12405 26 25 12439 SDFFRXL $T=1235100 1259110 0 0 $X=1235098 $Y=1258858
X446 11396 12389 12365 10868 9644 12221 26 25 12216 SDFFRXL $T=1246140 1251730 0 180 $X=1235100 $Y=1247790
X447 11737 11942 12250 10868 9644 10777 26 25 12445 SDFFRXL $T=1235560 1288630 1 0 $X=1235558 $Y=1284690
X448 12313 12379 12378 11826 11850 12237 26 25 12211 SDFFRXL $T=1246600 1192690 0 180 $X=1235560 $Y=1188750
X449 12452 12330 235 10868 9644 12259 26 25 12250 SDFFRXL $T=1248900 1281250 1 180 $X=1237860 $Y=1280998
X450 11396 12420 12439 10868 9644 12581 26 25 12642 SDFFRXL $T=1244760 1266490 0 0 $X=1244758 $Y=1266238
X451 233 248 247 243 99 12349 26 25 162 SDFFRXL $T=1256260 1347670 1 180 $X=1245220 $Y=1347418
X452 11396 236 12170 11826 11426 12693 26 25 12598 SDFFRXL $T=1247520 1229590 0 0 $X=1247518 $Y=1229338
X453 11396 12694 12676 10868 11850 12468 26 25 12195 SDFFRXL $T=1259020 1259110 1 180 $X=1247980 $Y=1258858
X454 12313 12767 258 11826 11850 12378 26 25 12565 SDFFRXL $T=1262700 1192690 0 180 $X=1251660 $Y=1188750
X455 12452 244 12606 10868 11270 12817 26 25 12747 SDFFRXL $T=1252580 1281250 0 0 $X=1252578 $Y=1280998
X456 12313 12781 12776 11826 9557 12596 26 25 12365 SDFFRXL $T=1263620 1200070 0 180 $X=1252580 $Y=1196130
X457 12452 12803 12677 12746 11850 12606 26 25 12135 SDFFRXL $T=1263620 1273870 1 180 $X=1252580 $Y=1273618
X458 11396 246 12468 10868 11426 12828 26 25 12640 SDFFRXL $T=1253040 1259110 1 0 $X=1253038 $Y=1255170
X459 12452 265 12828 12746 11270 12677 26 25 12652 SDFFRXL $T=1266840 1266490 1 180 $X=1255800 $Y=1266238
X460 233 12835 263 243 99 251 26 25 12626 SDFFRXL $T=1267300 1347670 1 180 $X=1256260 $Y=1347418
X461 12313 13008 12895 11826 9557 11335 26 25 12796 SDFFRXL $T=1273280 1185310 0 180 $X=1262240 $Y=1181370
X462 11396 12858 12852 12746 11850 13080 26 25 12238 SDFFRXL $T=1265000 1259110 1 0 $X=1264998 $Y=1255170
X463 11396 13066 12983 11826 11850 12852 26 25 12580 SDFFRXL $T=1276040 1236970 0 180 $X=1265000 $Y=1233030
X464 13081 13024 12817 12746 99 12859 26 25 11484 SDFFRXL $T=1276040 1296010 1 180 $X=1265000 $Y=1295758
X465 13081 13025 12859 12746 99 267 26 25 12215 SDFFRXL $T=1276040 1303390 1 180 $X=1265000 $Y=1303138
X466 12313 12911 12928 11826 9557 12867 26 25 13145 SDFFRXL $T=1266840 1185310 0 0 $X=1266838 $Y=1185058
X467 12452 12986 13080 12746 11850 12676 26 25 12503 SDFFRXL $T=1277880 1266490 0 180 $X=1266840 $Y=1262550
X468 12313 12896 13093 11826 9557 12876 26 25 12895 SDFFRXL $T=1278340 1192690 1 180 $X=1267300 $Y=1192438
X469 12313 12930 13094 11826 9815 12877 26 25 12897 SDFFRXL $T=1278340 1214830 0 180 $X=1267300 $Y=1210890
X470 12313 12945 13145 11826 9557 12962 26 25 12776 SDFFRXL $T=1280640 1200070 0 180 $X=1269600 $Y=1196130
X471 12313 12993 13009 11826 9815 13043 26 25 13094 SDFFRXL $T=1270060 1207450 0 0 $X=1270058 $Y=1207198
X472 11396 13183 12693 11826 11850 12983 26 25 12335 SDFFRXL $T=1281100 1229590 1 180 $X=1270060 $Y=1229338
X473 12313 13102 288 11826 9815 13032 26 25 13009 SDFFRXL $T=1283860 1200070 1 180 $X=1272820 $Y=1199818
X474 12313 13237 284 11826 9557 13056 26 25 12928 SDFFRXL $T=1284320 1185310 0 180 $X=1273280 $Y=1181370
X475 13081 13229 13260 243 147 13437 26 25 290 SDFFRXL $T=1282480 1347670 1 0 $X=1282478 $Y=1343730
X476 12313 13272 12897 11826 11426 13439 26 25 13273 SDFFRXL $T=1283860 1214830 1 0 $X=1283858 $Y=1210890
X477 11396 13313 13338 11826 147 13457 26 25 13380 SDFFRXL $T=1285700 1236970 1 0 $X=1285698 $Y=1233030
X478 13081 324 322 243 318 13316 26 25 303 SDFFRXL $T=1296740 1347670 1 180 $X=1285700 $Y=1347418
X479 12313 13348 13273 11826 11426 13513 26 25 13379 SDFFRXL $T=1287080 1214830 0 0 $X=1287078 $Y=1214578
X480 12313 13327 13257 11826 11426 13512 26 25 13256 SDFFRXL $T=1287540 1207450 1 0 $X=1287538 $Y=1203510
X481 12313 13328 13379 11826 11426 13511 26 25 13257 SDFFRXL $T=1287540 1207450 0 0 $X=1287538 $Y=1207198
X482 13349 13364 13380 12746 306 13476 26 25 13505 SDFFRXL $T=1287540 1251730 0 0 $X=1287538 $Y=1251478
X483 13081 13514 13382 12746 147 13366 26 25 13260 SDFFRXL $T=1298580 1325530 1 180 $X=1287540 $Y=1325278
X484 12452 13339 13388 12746 306 13548 26 25 13314 SDFFRXL $T=1288000 1266490 1 0 $X=1287998 $Y=1262550
X485 12313 13503 13502 11826 11426 13373 26 25 13093 SDFFRXL $T=1299040 1192690 1 180 $X=1288000 $Y=1192438
X486 13081 13352 310 12746 147 13559 26 25 13315 SDFFRXL $T=1288920 1340290 1 0 $X=1288918 $Y=1336350
X487 13081 13585 13445 12746 147 13430 26 25 13351 SDFFRXL $T=1301800 1296010 1 180 $X=1290760 $Y=1295758
X488 13349 13530 13458 11826 147 13590 26 25 13338 SDFFRXL $T=1296740 1236970 1 0 $X=1296738 $Y=1233030
X489 13081 13653 13693 12746 147 13616 26 25 13603 SDFFRXL $T=1312380 1318150 1 180 $X=1301340 $Y=1317898
X490 12313 13644 13663 11826 11426 13729 26 25 13608 SDFFRXL $T=1303180 1207450 0 0 $X=1303178 $Y=1207198
X491 15941 16427 16349 595 16449 16496 26 25 16490 SDFFRXL $T=1564460 1310770 0 0 $X=1564458 $Y=1310518
X492 15941 16428 16439 595 9816 16482 26 25 16491 SDFFRXL $T=1564460 1347670 1 0 $X=1564458 $Y=1343730
X493 15942 16434 16441 16011 16449 16421 26 25 16551 SDFFRXL $T=1564920 1281250 0 0 $X=1564918 $Y=1280998
X494 16334 16514 16495 16011 16483 16438 26 25 16432 SDFFRXL $T=1576420 1229590 1 180 $X=1565380 $Y=1229338
X495 16334 16518 16340 16011 16449 16413 26 25 16435 SDFFRXL $T=1576880 1259110 0 180 $X=1565840 $Y=1255170
X496 15937 16453 16466 16011 16483 16495 26 25 16566 SDFFRXL $T=1568600 1222210 0 0 $X=1568598 $Y=1221958
X497 610 16548 16541 595 9816 16439 26 25 16526 SDFFRXL $T=1587460 1340290 1 180 $X=1576420 $Y=1340038
X498 16334 16538 16438 16011 16483 16542 26 25 16622 SDFFRXL $T=1576880 1236970 1 0 $X=1576878 $Y=1233030
X499 16334 16525 16542 16011 16449 16510 26 25 16623 SDFFRXL $T=1576880 1244350 1 0 $X=1576878 $Y=1240410
X500 16334 16539 16510 16011 16449 16581 26 25 16616 SDFFRXL $T=1576880 1251730 1 0 $X=1576878 $Y=1247790
X501 15941 16540 16543 595 16449 16552 26 25 16617 SDFFRXL $T=1576880 1296010 0 0 $X=1576878 $Y=1295758
X502 15942 16605 16600 16011 16449 16362 26 25 16530 SDFFRXL $T=1587920 1266490 1 180 $X=1576880 $Y=1266238
X503 16334 16515 16412 16011 16449 16444 26 25 16631 SDFFRXL $T=1577340 1244350 0 0 $X=1577338 $Y=1244098
X504 16567 16598 16552 595 16449 16541 26 25 16533 SDFFRXL $T=1588380 1310770 0 180 $X=1577340 $Y=1306830
X505 15941 16529 16602 595 9816 16486 26 25 16534 SDFFRXL $T=1588380 1325530 1 180 $X=1577340 $Y=1325278
X506 15942 16547 16546 595 16449 16543 26 25 16553 SDFFRXL $T=1590680 1296010 0 180 $X=1579640 $Y=1292070
X507 610 16624 16620 595 76 16554 26 25 16544 SDFFRXL $T=1590680 1347670 0 180 $X=1579640 $Y=1343730
X508 16567 16582 16421 16011 16483 16627 26 25 16635 SDFFRXL $T=1581020 1281250 0 0 $X=1581018 $Y=1280998
X509 16567 16563 16581 16011 16483 16545 26 25 16633 SDFFRXL $T=1581480 1266490 1 0 $X=1581478 $Y=1262550
X510 16567 16564 16545 16011 16449 16546 26 25 16621 SDFFRXL $T=1581480 1273870 1 0 $X=1581478 $Y=1269930
X511 15941 16588 16568 595 9816 16602 26 25 16675 SDFFRXL $T=1581940 1310770 0 0 $X=1581938 $Y=1310518
X512 562 16589 608 595 76 16620 26 25 16634 SDFFRXL $T=1581940 1347670 0 0 $X=1581938 $Y=1347418
X513 16334 16612 16626 16011 16483 16466 26 25 16583 SDFFRXL $T=1592980 1222210 1 180 $X=1581940 $Y=1221958
X514 15941 16593 16594 595 9816 16568 26 25 16696 SDFFRXL $T=1582400 1325530 1 0 $X=1582398 $Y=1321590
X515 610 16632 16646 595 9816 16594 26 25 16586 SDFFRXL $T=1593440 1332910 1 180 $X=1582400 $Y=1332658
X516 16567 16723 16719 595 16483 16645 26 25 16629 SDFFRXL $T=1601720 1296010 0 180 $X=1590680 $Y=1292070
X517 16567 16673 16683 16011 16483 16693 26 25 16761 SDFFRXL $T=1591600 1273870 0 0 $X=1591598 $Y=1273618
X518 16567 16674 16684 595 16483 16719 26 25 16764 SDFFRXL $T=1591600 1303390 0 0 $X=1591598 $Y=1303138
X519 16567 16711 16762 595 9816 16684 26 25 16679 SDFFRXL $T=1604020 1310770 1 180 $X=1592980 $Y=1310518
X520 16334 16690 16692 16011 16483 16765 26 25 16780 SDFFRXL $T=1593440 1251730 1 0 $X=1593438 $Y=1247790
X521 16567 16766 16645 16011 16483 16688 26 25 16651 SDFFRXL $T=1604480 1288630 0 180 $X=1593440 $Y=1284690
X522 16567 16691 16702 16011 16483 16692 26 25 16786 SDFFRXL $T=1594820 1259110 1 0 $X=1594818 $Y=1255170
X523 610 16697 16703 595 9816 16646 26 25 16773 SDFFRXL $T=1594820 1332910 0 0 $X=1594818 $Y=1332658
X524 16567 16770 16627 16011 16483 16683 26 25 16650 SDFFRXL $T=1606320 1281250 0 180 $X=1595280 $Y=1277310
X525 16334 16771 16714 16011 16483 16626 26 25 16698 SDFFRXL $T=1606780 1222210 1 180 $X=1595740 $Y=1221958
X526 16334 16775 16765 16011 16483 16714 26 25 16710 SDFFRXL $T=1608160 1236970 0 180 $X=1597120 $Y=1233030
X527 610 627 16554 595 622 620 26 25 16654 SDFFRXL $T=1609080 1347670 0 180 $X=1598040 $Y=1343730
X528 16567 16731 16693 16011 16483 16600 26 25 16781 SDFFRXL $T=1598960 1273870 1 0 $X=1598958 $Y=1269930
X529 16567 16732 16688 16011 16483 16783 26 25 16787 SDFFRXL $T=1598960 1288630 0 0 $X=1598958 $Y=1288378
X530 610 16733 323 595 9816 16703 26 25 16772 SDFFRXL $T=1598960 1332910 1 0 $X=1598958 $Y=1328970
X531 16567 16769 16778 16011 16483 16702 26 25 16724 SDFFRXL $T=1610000 1259110 1 180 $X=1598960 $Y=1258858
X532 16567 16819 16783 595 16449 16763 26 25 16648 SDFFRXL $T=1612760 1296010 0 180 $X=1601720 $Y=1292070
X533 16567 16822 16763 16011 16483 16767 26 25 16653 SDFFRXL $T=1613680 1273870 1 180 $X=1602640 $Y=1273618
X534 16567 16821 16820 595 16449 16768 26 25 16613 SDFFRXL $T=1613680 1303390 1 180 $X=1602640 $Y=1303138
X535 16567 16826 16768 595 16449 16762 26 25 16652 SDFFRXL $T=1615060 1310770 1 180 $X=1604020 $Y=1310518
X536 16567 16830 16767 16011 16483 16778 26 25 16628 SDFFRXL $T=1621960 1266490 1 180 $X=1610920 $Y=1266238
X537 610 16847 16831 595 622 16823 26 25 16716 SDFFRXL $T=1622880 1325530 1 180 $X=1611840 $Y=1325278
X538 610 16848 630 595 622 16824 26 25 16725 SDFFRXL $T=1622880 1347670 0 180 $X=1611840 $Y=1343730
X539 16567 16879 16834 595 16449 16820 26 25 16516 SDFFRXL $T=1623340 1303390 0 180 $X=1612300 $Y=1299450
X540 610 636 633 595 622 630 26 25 16782 SDFFRXL $T=1623340 1347670 1 180 $X=1612300 $Y=1347418
X541 610 16829 16832 595 622 16831 26 25 16595 SDFFRXL $T=1625640 1332910 0 180 $X=1614600 $Y=1328970
X542 610 16880 16824 595 622 16832 26 25 16779 SDFFRXL $T=1625640 1340290 1 180 $X=1614600 $Y=1340038
X543 610 16886 16823 595 622 16834 26 25 16712 SDFFRXL $T=1626100 1325530 0 180 $X=1615060 $Y=1321590
X544 8948 25 8951 26 CLKBUFX2 $T=1065820 1192690 0 0 $X=1065818 $Y=1192438
X545 32 25 9557 26 CLKBUFX2 $T=1104920 1303390 0 0 $X=1104918 $Y=1303138
X546 9664 25 9069 26 CLKBUFX2 $T=1109060 1325530 1 0 $X=1109058 $Y=1321590
X547 9705 25 68 26 CLKBUFX2 $T=1110900 1325530 1 0 $X=1110898 $Y=1321590
X548 66 25 9547 26 CLKBUFX2 $T=1112740 1318150 1 180 $X=1110900 $Y=1317898
X549 85 25 9382 26 CLKBUFX2 $T=1121020 1266490 0 0 $X=1121018 $Y=1266238
X550 9776 25 91 26 CLKBUFX2 $T=1121020 1347670 1 0 $X=1121018 $Y=1343730
X551 89 25 9723 26 CLKBUFX2 $T=1123320 1325530 1 180 $X=1121480 $Y=1325278
X552 44 25 9963 26 CLKBUFX2 $T=1121940 1236970 0 0 $X=1121938 $Y=1236718
X553 9931 25 71 26 CLKBUFX2 $T=1122860 1332910 0 0 $X=1122858 $Y=1332658
X554 96 25 9930 26 CLKBUFX2 $T=1128380 1332910 1 180 $X=1126540 $Y=1332658
X555 10104 25 69 26 CLKBUFX2 $T=1129760 1340290 0 0 $X=1129758 $Y=1340038
X556 10147 25 10122 26 CLKBUFX2 $T=1131140 1266490 1 0 $X=1131138 $Y=1262550
X557 9570 25 10216 26 CLKBUFX2 $T=1132520 1148410 1 0 $X=1132518 $Y=1144470
X558 9393 25 10176 26 CLKBUFX2 $T=1134820 1133650 1 0 $X=1134818 $Y=1129710
X559 10209 25 10260 26 CLKBUFX2 $T=1135280 1288630 1 0 $X=1135278 $Y=1284690
X560 9686 25 10273 26 CLKBUFX2 $T=1136660 1207450 1 0 $X=1136658 $Y=1203510
X561 10281 25 10290 26 CLKBUFX2 $T=1139420 1288630 1 0 $X=1139418 $Y=1284690
X562 9897 25 10373 26 CLKBUFX2 $T=1140800 1207450 0 0 $X=1140798 $Y=1207198
X563 9740 25 10417 26 CLKBUFX2 $T=1141260 1148410 1 0 $X=1141258 $Y=1144470
X564 10362 25 10045 26 CLKBUFX2 $T=1141260 1281250 1 0 $X=1141258 $Y=1277310
X565 10322 25 10331 26 CLKBUFX2 $T=1145400 1111510 1 0 $X=1145398 $Y=1107570
X566 10004 25 10191 26 CLKBUFX2 $T=1153220 1259110 0 0 $X=1153218 $Y=1258858
X567 9525 25 10807 26 CLKBUFX2 $T=1163340 1177930 0 0 $X=1163338 $Y=1177678
X568 10599 25 9664 26 CLKBUFX2 $T=1163340 1310770 0 0 $X=1163338 $Y=1310518
X569 10755 25 10055 26 CLKBUFX2 $T=1163800 1074610 0 0 $X=1163798 $Y=1074358
X570 10869 25 10067 26 CLKBUFX2 $T=1168860 1273870 0 0 $X=1168858 $Y=1273618
X571 10472 25 10972 26 CLKBUFX2 $T=1170240 1222210 0 0 $X=1170238 $Y=1221958
X572 10750 25 10935 26 CLKBUFX2 $T=1171160 1052470 0 0 $X=1171158 $Y=1052218
X573 10887 25 9916 26 CLKBUFX2 $T=1173920 1104130 1 0 $X=1173918 $Y=1100190
X574 10521 25 9780 26 CLKBUFX2 $T=1176220 1222210 0 0 $X=1176218 $Y=1221958
X575 10908 25 11242 26 CLKBUFX2 $T=1186340 1133650 0 0 $X=1186338 $Y=1133398
X576 10290 25 10426 26 CLKBUFX2 $T=1188640 1251730 1 0 $X=1188638 $Y=1247790
X577 10750 25 10764 26 CLKBUFX2 $T=1193240 1148410 1 0 $X=1193238 $Y=1144470
X578 11396 25 10521 26 CLKBUFX2 $T=1199680 1236970 1 0 $X=1199678 $Y=1233030
X579 11206 25 11241 26 CLKBUFX2 $T=1210260 1037710 1 0 $X=1210258 $Y=1033770
X580 11737 25 10599 26 CLKBUFX2 $T=1214400 1296010 0 0 $X=1214398 $Y=1295758
X581 11780 25 11821 26 CLKBUFX2 $T=1214860 1273870 0 0 $X=1214858 $Y=1273618
X582 12016 25 12005 26 CLKBUFX2 $T=1226820 1273870 1 0 $X=1226818 $Y=1269930
X583 12015 25 12017 26 CLKBUFX2 $T=1228660 1259110 1 0 $X=1228658 $Y=1255170
X584 10417 25 12364 26 CLKBUFX2 $T=1239700 1148410 1 0 $X=1239698 $Y=1144470
X585 12336 25 12000 26 CLKBUFX2 $T=1242460 1325530 1 0 $X=1242458 $Y=1321590
X586 12117 25 12001 26 CLKBUFX2 $T=1257640 1325530 1 0 $X=1257638 $Y=1321590
X587 12452 25 11396 26 CLKBUFX2 $T=1265000 1266490 1 0 $X=1264998 $Y=1262550
X588 13032 25 13233 26 CLKBUFX2 $T=1278340 1222210 1 0 $X=1278338 $Y=1218270
X589 12867 25 13227 26 CLKBUFX2 $T=1279260 1185310 0 0 $X=1279258 $Y=1185058
X590 12962 25 13293 26 CLKBUFX2 $T=1282480 1236970 0 0 $X=1282478 $Y=1236718
X591 13056 25 13387 26 CLKBUFX2 $T=1288000 1177930 0 0 $X=1287998 $Y=1177678
X592 201 25 11270 26 CLKBUFX2 $T=1290760 1318150 1 0 $X=1290758 $Y=1314210
X593 13043 25 13563 26 CLKBUFX2 $T=1294440 1222210 1 0 $X=1294438 $Y=1218270
X594 13609 25 12313 26 CLKBUFX2 $T=1301340 1207450 0 0 $X=1301338 $Y=1207198
X595 13646 25 13349 26 CLKBUFX2 $T=1303180 1251730 0 0 $X=1303178 $Y=1251478
X596 13349 25 13609 26 CLKBUFX2 $T=1307320 1222210 1 0 $X=1307318 $Y=1218270
X597 13640 25 13560 26 CLKBUFX2 $T=1315140 1141030 1 0 $X=1315138 $Y=1137090
X598 348 25 13081 26 CLKBUFX2 $T=1315140 1332910 0 0 $X=1315138 $Y=1332658
X599 348 25 392 26 CLKBUFX2 $T=1337220 1347670 1 0 $X=1337218 $Y=1343730
X600 12452 25 13566 26 CLKBUFX2 $T=1338140 1296010 1 0 $X=1338138 $Y=1292070
X601 397 25 13851 26 CLKBUFX2 $T=1346420 1340290 1 0 $X=1346418 $Y=1336350
X602 14284 25 13640 26 CLKBUFX2 $T=1366200 1104130 1 0 $X=1366198 $Y=1100190
X603 14732 25 14465 26 CLKBUFX2 $T=1401160 1222210 1 0 $X=1401158 $Y=1218270
X604 14518 25 14400 26 CLKBUFX2 $T=1402540 1133650 1 0 $X=1402538 $Y=1129710
X605 14639 25 463 26 CLKBUFX2 $T=1403920 1340290 0 0 $X=1403918 $Y=1340038
X606 466 25 14596 26 CLKBUFX2 $T=1406680 1347670 0 0 $X=1406678 $Y=1347418
X607 459 25 14673 26 CLKBUFX2 $T=1412660 1347670 1 0 $X=1412658 $Y=1343730
X608 362 25 477 26 CLKBUFX2 $T=1418640 1340290 0 0 $X=1418638 $Y=1340038
X609 14751 25 14607 26 CLKBUFX2 $T=1422320 1259110 1 0 $X=1422318 $Y=1255170
X610 474 25 14773 26 CLKBUFX2 $T=1423700 1347670 1 0 $X=1423698 $Y=1343730
X611 484 25 14599 26 CLKBUFX2 $T=1425540 1347670 1 0 $X=1425538 $Y=1343730
X612 15135 25 14751 26 CLKBUFX2 $T=1452220 1236970 1 0 $X=1452218 $Y=1233030
X613 15292 25 14150 26 CLKBUFX2 $T=1459120 1281250 0 0 $X=1459118 $Y=1280998
X614 15353 25 14284 26 CLKBUFX2 $T=1466480 1126270 1 0 $X=1466478 $Y=1122330
X615 14868 25 15358 26 CLKBUFX2 $T=1468780 1192690 1 0 $X=1468778 $Y=1188750
X616 15353 25 14868 26 CLKBUFX2 $T=1472000 1207450 1 0 $X=1471998 $Y=1203510
X617 494 25 15225 26 CLKBUFX2 $T=1472000 1347670 0 0 $X=1471998 $Y=1347418
X618 15437 25 15135 26 CLKBUFX2 $T=1474760 1259110 1 0 $X=1474758 $Y=1255170
X619 15358 25 15293 26 CLKBUFX2 $T=1477060 1163170 1 0 $X=1477058 $Y=1159230
X620 513 25 15247 26 CLKBUFX2 $T=1508800 1325530 1 0 $X=1508798 $Y=1321590
X621 15760 25 15292 26 CLKBUFX2 $T=1515240 1296010 1 0 $X=1515238 $Y=1292070
X622 549 25 15321 26 CLKBUFX2 $T=1515700 1325530 0 0 $X=1515698 $Y=1325278
X623 90 25 550 26 CLKBUFX2 $T=1519840 1347670 1 0 $X=1519838 $Y=1343730
X624 555 25 15692 26 CLKBUFX2 $T=1523980 1273870 0 0 $X=1523978 $Y=1273618
X625 15631 25 14732 26 CLKBUFX2 $T=1524900 1229590 0 0 $X=1524898 $Y=1229338
X626 568 25 16189 26 CLKBUFX2 $T=1543300 1347670 0 0 $X=1543298 $Y=1347418
X627 536 25 577 26 CLKBUFX2 $T=1545140 1347670 0 0 $X=1545138 $Y=1347418
X628 15996 25 589 26 CLKBUFX2 $T=1552500 1347670 0 0 $X=1552498 $Y=1347418
X629 15937 25 15926 26 CLKBUFX2 $T=1560780 1192690 0 0 $X=1560778 $Y=1192438
X630 15942 25 16334 26 CLKBUFX2 $T=1569980 1266490 0 0 $X=1569978 $Y=1266238
X631 16486 25 598 26 CLKBUFX2 $T=1573200 1332910 0 180 $X=1571360 $Y=1328970
X632 16334 25 15937 26 CLKBUFX2 $T=1575500 1222210 1 0 $X=1575498 $Y=1218270
X633 15941 25 16567 26 CLKBUFX2 $T=1580100 1310770 0 0 $X=1580098 $Y=1310518
X634 603 25 16519 26 CLKBUFX2 $T=1585160 1318150 1 0 $X=1585158 $Y=1314210
X635 610 25 15941 26 CLKBUFX2 $T=1586540 1332910 1 0 $X=1586538 $Y=1328970
X636 16485 25 16442 26 CLKBUFX2 $T=1593900 1296010 0 0 $X=1593898 $Y=1295758
X637 129 25 13726 26 CLKBUFX2 $T=1595280 1340290 0 0 $X=1595278 $Y=1340038
X638 604 25 16414 26 CLKBUFX2 $T=1598960 1296010 0 0 $X=1598958 $Y=1295758
X639 625 25 16485 26 CLKBUFX2 $T=1606780 1332910 0 0 $X=1606778 $Y=1332658
X640 16449 25 16483 26 CLKBUFX2 $T=1612760 1296010 1 0 $X=1612758 $Y=1292070
X641 16825 25 16400 26 CLKBUFX2 $T=1614140 1310770 1 0 $X=1614138 $Y=1306830
X642 619 25 16825 26 CLKBUFX2 $T=1615980 1340290 1 0 $X=1615978 $Y=1336350
X643 9428 9619 9416 25 26 9546 MX2XL $T=1107220 1229590 0 180 $X=1103540 $Y=1225650
X644 67 69 28 25 26 9669 MX2XL $T=1113200 1340290 1 180 $X=1109520 $Y=1340038
X645 9678 9689 9735 25 26 9811 MX2XL $T=1109980 1133650 0 0 $X=1109978 $Y=1133398
X646 67 71 31 25 26 9682 MX2XL $T=1113660 1332910 1 180 $X=1109980 $Y=1332658
X647 67 68 9419 25 26 9783 MX2XL $T=1111820 1325530 0 0 $X=1111818 $Y=1325278
X648 9779 9797 9847 25 26 9910 MX2XL $T=1115500 1111510 0 0 $X=1115498 $Y=1111258
X649 9680 9813 9870 25 26 9896 MX2XL $T=1116880 1192690 0 0 $X=1116878 $Y=1192438
X650 9812 9859 9912 25 26 10029 MX2XL $T=1119180 1170550 1 0 $X=1119178 $Y=1166610
X651 9884 9875 9947 25 26 10038 MX2XL $T=1120560 1118890 0 0 $X=1120558 $Y=1118638
X652 9836 9798 9961 25 26 9990 MX2XL $T=1121020 1148410 0 0 $X=1121018 $Y=1148158
X653 67 91 57 25 26 9977 MX2XL $T=1129300 1347670 0 180 $X=1125620 $Y=1343730
X654 9170 10030 10101 25 26 10183 MX2XL $T=1127460 1177930 0 0 $X=1127458 $Y=1177678
X655 10055 8736 8732 25 26 10246 MX2XL $T=1128380 1074610 1 0 $X=1128378 $Y=1070670
X656 10055 8732 8742 25 26 10151 MX2XL $T=1128380 1074610 0 0 $X=1128378 $Y=1074358
X657 10057 9989 10137 25 26 10119 MX2XL $T=1128380 1148410 1 0 $X=1128378 $Y=1144470
X658 10061 10097 10155 25 26 10268 MX2XL $T=1129300 1163170 1 0 $X=1129298 $Y=1159230
X659 10055 8871 8736 25 26 10221 MX2XL $T=1131140 1089370 0 0 $X=1131138 $Y=1089118
X660 10055 8883 8871 25 26 10255 MX2XL $T=1131600 1081990 0 0 $X=1131598 $Y=1081738
X661 10055 8814 8816 25 26 10387 MX2XL $T=1132060 1067230 1 0 $X=1132058 $Y=1063290
X662 10055 8742 8748 25 26 10308 MX2XL $T=1136660 1067230 0 0 $X=1136658 $Y=1066978
X663 10211 10197 10295 25 26 10434 MX2XL $T=1136660 1133650 1 0 $X=1136658 $Y=1129710
X664 10055 8816 8749 25 26 10414 MX2XL $T=1144020 1074610 1 0 $X=1144018 $Y=1070670
X665 10332 10411 10479 25 26 10478 MX2XL $T=1144940 1141030 0 0 $X=1144938 $Y=1140778
X666 10055 8749 8961 25 26 10489 MX2XL $T=1145860 1059850 0 0 $X=1145858 $Y=1059598
X667 10055 8748 8814 25 26 10309 MX2XL $T=1153680 1074610 1 180 $X=1150000 $Y=1074358
X668 10055 9003 9101 25 26 10628 MX2XL $T=1154600 1059850 0 0 $X=1154598 $Y=1059598
X669 10055 8961 9003 25 26 10574 MX2XL $T=1159660 1074610 0 180 $X=1155980 $Y=1070670
X670 10055 9270 9386 25 26 10786 MX2XL $T=1161040 1059850 0 0 $X=1161038 $Y=1059598
X671 10055 9101 9228 25 26 10671 MX2XL $T=1165180 1074610 0 180 $X=1161500 $Y=1070670
X672 10750 9101 9003 25 26 10916 MX2XL $T=1162880 1052470 1 0 $X=1162878 $Y=1048530
X673 10055 9228 9102 25 26 10603 MX2XL $T=1166560 1067230 0 180 $X=1162880 $Y=1063290
X674 10755 9102 9270 25 26 10793 MX2XL $T=1163340 1081990 0 0 $X=1163338 $Y=1081738
X675 10750 9003 8961 25 26 10883 MX2XL $T=1165180 1059850 0 0 $X=1165178 $Y=1059598
X676 10750 8816 8814 25 26 10903 MX2XL $T=1167020 1059850 1 0 $X=1167018 $Y=1055910
X677 10750 8961 8749 25 26 10915 MX2XL $T=1167480 1045090 0 0 $X=1167478 $Y=1044838
X678 10470 8742 8732 25 26 10928 MX2XL $T=1167480 1074610 1 0 $X=1167478 $Y=1070670
X679 10750 8749 8816 25 26 10944 MX2XL $T=1169780 1059850 0 0 $X=1169778 $Y=1059598
X680 10750 9102 9228 25 26 11078 MX2XL $T=1171620 1052470 1 0 $X=1171618 $Y=1048530
X681 10750 8748 8742 25 26 10965 MX2XL $T=1171620 1067230 1 0 $X=1171618 $Y=1063290
X682 10750 8814 8748 25 26 11039 MX2XL $T=1171620 1067230 0 0 $X=1171618 $Y=1066978
X683 10750 9228 9101 25 26 11106 MX2XL $T=1173000 1059850 1 0 $X=1172998 $Y=1055910
X684 10750 8732 8736 25 26 11004 MX2XL $T=1173000 1074610 1 0 $X=1172998 $Y=1070670
X685 10755 9386 11066 25 26 10745 MX2XL $T=1182200 1081990 1 180 $X=1178520 $Y=1081738
X686 10755 11063 11087 25 26 10852 MX2XL $T=1183120 1096750 0 180 $X=1179440 $Y=1092810
X687 10935 9270 9102 25 26 11105 MX2XL $T=1184040 1052470 1 180 $X=1180360 $Y=1052218
X688 10755 11066 11063 25 26 10890 MX2XL $T=1184500 1081990 0 180 $X=1180820 $Y=1078050
X689 10750 8871 8883 25 26 11160 MX2XL $T=1181280 1074610 0 0 $X=1181278 $Y=1074358
X690 10755 11087 11225 25 26 10936 MX2XL $T=1184500 1081990 0 0 $X=1184498 $Y=1081738
X691 10935 11066 9386 25 26 11379 MX2XL $T=1188640 1059850 1 0 $X=1188638 $Y=1055910
X692 10935 9386 9270 25 26 11268 MX2XL $T=1192780 1052470 1 180 $X=1189100 $Y=1052218
X693 10755 10967 11052 25 26 11280 MX2XL $T=1193700 1104130 0 180 $X=1190020 $Y=1100190
X694 10755 11225 11244 25 26 11080 MX2XL $T=1193700 1111510 0 180 $X=1190020 $Y=1107570
X695 10755 11244 11295 25 26 11258 MX2XL $T=1194160 1081990 1 180 $X=1190480 $Y=1081738
X696 10755 11323 11023 25 26 11320 MX2XL $T=1200140 1096750 1 180 $X=1196460 $Y=1096498
X697 10755 11344 11275 25 26 11259 MX2XL $T=1200140 1111510 1 180 $X=1196460 $Y=1111258
X698 10755 11243 11344 25 26 11331 MX2XL $T=1200600 1089370 1 180 $X=1196920 $Y=1089118
X699 10755 11147 11437 25 26 11279 MX2XL $T=1201520 1104130 0 180 $X=1197840 $Y=1100190
X700 10755 11295 11243 25 26 11171 MX2XL $T=1201520 1111510 0 180 $X=1197840 $Y=1107570
X701 10755 11275 11322 25 26 11284 MX2XL $T=1201980 1096750 0 180 $X=1198300 $Y=1092810
X702 10935 11063 11066 25 26 11629 MX2XL $T=1208420 1059850 1 0 $X=1208418 $Y=1055910
X703 10935 11052 10967 25 26 11838 MX2XL $T=1214860 1089370 0 0 $X=1214858 $Y=1089118
X704 10935 11087 11063 25 26 11724 MX2XL $T=1221760 1059850 1 180 $X=1218080 $Y=1059598
X705 10935 10967 11437 25 26 11797 MX2XL $T=1223140 1096750 0 180 $X=1219460 $Y=1092810
X706 10935 11147 11023 25 26 11933 MX2XL $T=1227280 1089370 1 180 $X=1223600 $Y=1089118
X707 10935 11323 11322 25 26 12012 MX2XL $T=1224980 1089370 1 0 $X=1224978 $Y=1085430
X708 10935 11275 11344 25 26 12003 MX2XL $T=1234640 1081990 1 180 $X=1230960 $Y=1081738
X709 10935 11437 11147 25 26 12053 MX2XL $T=1234640 1089370 1 180 $X=1230960 $Y=1089118
X710 10935 11344 11243 25 26 12113 MX2XL $T=1231420 1081990 1 0 $X=1231418 $Y=1078050
X711 10935 11295 11244 25 26 12126 MX2XL $T=1236480 1074610 0 180 $X=1232800 $Y=1070670
X712 10935 11243 11295 25 26 12054 MX2XL $T=1236480 1074610 1 180 $X=1232800 $Y=1074358
X713 10935 11225 11087 25 26 11847 MX2XL $T=1239700 1067230 0 180 $X=1236020 $Y=1063290
X714 10935 11244 11225 25 26 11794 MX2XL $T=1241080 1067230 1 180 $X=1237400 $Y=1066978
X715 10935 11322 11275 25 26 12222 MX2XL $T=1241080 1081990 1 180 $X=1237400 $Y=1081738
X716 10935 11023 11323 25 26 12174 MX2XL $T=1241080 1089370 1 180 $X=1237400 $Y=1089118
X717 586 13235 581 25 26 16198 MX2XL $T=1550660 1340290 0 180 $X=1546980 $Y=1336350
X718 586 13679 582 25 26 579 MX2XL $T=1551120 1347670 1 180 $X=1547440 $Y=1347418
X719 586 14741 16215 25 26 16330 MX2XL $T=1553420 1332910 1 0 $X=1553418 $Y=1328970
X720 586 13843 16204 25 26 16315 MX2XL $T=1553880 1325530 1 0 $X=1553878 $Y=1321590
X721 587 13958 16390 25 26 16404 MX2XL $T=1558940 1200070 1 0 $X=1558938 $Y=1196130
X722 587 14833 16391 25 26 16405 MX2XL $T=1558940 1207450 1 0 $X=1558938 $Y=1203510
X723 587 14458 16369 25 26 16406 MX2XL $T=1558940 1214830 1 0 $X=1558938 $Y=1210890
X724 586 13725 16343 25 26 16398 MX2XL $T=1558940 1303390 1 0 $X=1558938 $Y=1299450
X725 587 13350 16349 25 26 16415 MX2XL $T=1559400 1310770 0 0 $X=1559398 $Y=1310518
X726 586 13629 16396 25 26 16371 MX2XL $T=1559400 1347670 1 0 $X=1559398 $Y=1343730
X727 587 13567 16358 25 26 16425 MX2XL $T=1561240 1229590 0 0 $X=1561238 $Y=1229338
X728 587 13739 16412 25 26 16422 MX2XL $T=1561240 1244350 0 0 $X=1561238 $Y=1244098
X729 586 13786 16332 25 26 16419 MX2XL $T=1561240 1340290 1 0 $X=1561238 $Y=1336350
X730 587 13971 16186 25 26 16328 MX2XL $T=1564920 1288630 1 180 $X=1561240 $Y=1288378
X731 586 13717 16399 25 26 16469 MX2XL $T=1561700 1332910 1 0 $X=1561698 $Y=1328970
X732 587 13919 16394 25 26 16503 MX2XL $T=1563540 1296010 1 0 $X=1563538 $Y=1292070
X733 587 14743 16340 25 26 16450 MX2XL $T=1565380 1251730 0 0 $X=1565378 $Y=1251478
X734 587 13471 16388 25 26 16456 MX2XL $T=1573200 1318150 1 180 $X=1569520 $Y=1317898
X735 587 14203 16310 25 26 16440 MX2XL $T=1573660 1229590 0 180 $X=1569980 $Y=1225650
X736 587 13689 16418 25 26 16484 MX2XL $T=1575500 1266490 1 180 $X=1571820 $Y=1266238
X737 587 13881 16468 25 26 16431 MX2XL $T=1586080 1214830 1 180 $X=1582400 $Y=1214578
X738 587 13782 16417 25 26 16504 MX2XL $T=1587000 1207450 1 180 $X=1583320 $Y=1207198
X739 587 13764 16368 25 26 16508 MX2XL $T=1591140 1192690 0 180 $X=1587460 $Y=1188750
X740 587 13902 16509 25 26 16430 MX2XL $T=1591140 1200070 1 180 $X=1587460 $Y=1199818
X741 10042 10331 10002 10399 25 26 MXI2X1 $T=1138960 1096750 1 0 $X=1138958 $Y=1092810
X742 10230 10322 10208 10389 25 26 MXI2X1 $T=1138960 1111510 0 0 $X=1138958 $Y=1111258
X743 10124 10331 10190 10493 25 26 MXI2X1 $T=1144480 1096750 1 0 $X=1144478 $Y=1092810
X744 10321 10331 10388 10490 25 26 MXI2X1 $T=1145860 1104130 0 0 $X=1145858 $Y=1103878
X745 10438 10322 10319 10538 25 26 MXI2X1 $T=1145860 1126270 1 0 $X=1145858 $Y=1122330
X746 10432 10266 10447 10241 25 26 MXI2X1 $T=1149080 1081990 1 180 $X=1145860 $Y=1081738
X747 10406 10331 10154 10526 25 26 MXI2X1 $T=1146320 1096750 0 0 $X=1146318 $Y=1096498
X748 10575 10266 10548 10463 25 26 MXI2X1 $T=1153680 1081990 0 180 $X=1150460 $Y=1078050
X749 10529 10266 10545 10257 25 26 MXI2X1 $T=1153680 1111510 1 180 $X=1150460 $Y=1111258
X750 10393 10322 10644 10615 25 26 MXI2X1 $T=1154600 1104130 0 0 $X=1154598 $Y=1103878
X751 10466 10322 10646 10709 25 26 MXI2X1 $T=1155520 1118890 0 0 $X=1155518 $Y=1118638
X752 10576 10207 10465 10675 25 26 MXI2X1 $T=1155980 1096750 1 0 $X=1155978 $Y=1092810
X753 10656 10266 10624 10529 25 26 MXI2X1 $T=1159200 1111510 1 180 $X=1155980 $Y=1111258
X754 10629 10207 10551 10684 25 26 MXI2X1 $T=1156440 1089370 1 0 $X=1156438 $Y=1085430
X755 10656 10207 10782 10763 25 26 MXI2X1 $T=1160580 1118890 0 0 $X=1160578 $Y=1118638
X756 10745 10185 10740 10793 25 26 MXI2X1 $T=1161960 1089370 0 0 $X=1161958 $Y=1089118
X757 10208 9916 10828 10866 25 26 MXI2X1 $T=1162420 1111510 0 0 $X=1162418 $Y=1111258
X758 10794 10266 10634 10740 25 26 MXI2X1 $T=1165640 1111510 0 180 $X=1162420 $Y=1107570
X759 10672 10207 10536 10929 25 26 MXI2X1 $T=1167480 1089370 0 0 $X=1167478 $Y=1089118
X760 10890 10185 10851 10786 25 26 MXI2X1 $T=1170700 1074610 1 180 $X=1167480 $Y=1074358
X761 10891 10266 10787 10851 25 26 MXI2X1 $T=1170700 1089370 0 180 $X=1167480 $Y=1085430
X762 10763 10207 10810 10922 25 26 MXI2X1 $T=1168860 1111510 0 0 $X=1168858 $Y=1111258
X763 10154 9916 10923 10904 25 26 MXI2X1 $T=1170240 1104130 1 0 $X=1170238 $Y=1100190
X764 10852 10299 10794 11080 25 26 MXI2X1 $T=1170700 1104130 0 0 $X=1170698 $Y=1103878
X765 10319 10887 11058 10921 25 26 MXI2X1 $T=1171620 1126270 1 0 $X=1171618 $Y=1122330
X766 10832 10871 10918 10811 25 26 MXI2X1 $T=1171620 1155790 0 0 $X=1171618 $Y=1155538
X767 10915 10951 10927 10903 25 26 MXI2X1 $T=1174840 1037710 0 180 $X=1171620 $Y=1033770
X768 10936 10185 10980 10890 25 26 MXI2X1 $T=1172080 1081990 0 0 $X=1172078 $Y=1081738
X769 10903 10951 11038 10965 25 26 MXI2X1 $T=1172540 1037710 0 0 $X=1172538 $Y=1037458
X770 10916 10951 10938 10915 25 26 MXI2X1 $T=1175760 1045090 0 180 $X=1172540 $Y=1041150
X771 10952 10266 10788 10980 25 26 MXI2X1 $T=1173000 1089370 0 0 $X=1172998 $Y=1089118
X772 10947 10871 11088 10901 25 26 MXI2X1 $T=1173460 1141030 1 0 $X=1173458 $Y=1137090
X773 10883 10951 10994 10944 25 26 MXI2X1 $T=1173920 1059850 0 0 $X=1173918 $Y=1059598
X774 11112 11133 10175 11061 25 26 MXI2X1 $T=1181740 1045090 0 180 $X=1178520 $Y=1041150
X775 11080 10299 11007 11171 25 26 MXI2X1 $T=1178980 1111510 1 0 $X=1178978 $Y=1107570
X776 10646 10887 11185 11094 25 26 MXI2X1 $T=1178980 1126270 1 0 $X=1178978 $Y=1122330
X777 10963 10871 11207 10756 25 26 MXI2X1 $T=1179440 1133650 0 0 $X=1179438 $Y=1133398
X778 11106 10951 11138 10883 25 26 MXI2X1 $T=1179900 1059850 0 0 $X=1179898 $Y=1059598
X779 10944 10951 11194 11039 25 26 MXI2X1 $T=1179900 1067230 1 0 $X=1179898 $Y=1063290
X780 10002 10887 11183 11093 25 26 MXI2X1 $T=1179900 1096750 0 0 $X=1179898 $Y=1096498
X781 10936 10299 10891 11258 25 26 MXI2X1 $T=1180360 1089370 1 0 $X=1180358 $Y=1085430
X782 11088 10605 11135 11172 25 26 MXI2X1 $T=1180360 1141030 1 0 $X=1180358 $Y=1137090
X783 11105 10951 11119 11106 25 26 MXI2X1 $T=1183580 1059850 0 180 $X=1180360 $Y=1055910
X784 10918 10908 10995 11083 25 26 MXI2X1 $T=1183580 1155790 1 180 $X=1180360 $Y=1155538
X785 11078 10951 11142 10916 25 26 MXI2X1 $T=1184960 1045090 1 180 $X=1181740 $Y=1044838
X786 11171 10299 10930 11259 25 26 MXI2X1 $T=1184500 1111510 1 0 $X=1184498 $Y=1107570
X787 11218 11133 10471 11272 25 26 MXI2X1 $T=1185880 1074610 0 0 $X=1185878 $Y=1074358
X788 11207 140 11260 11203 25 26 MXI2X1 $T=1185880 1141030 0 0 $X=1185878 $Y=1140778
X789 11259 10299 10962 11308 25 26 MXI2X1 $T=1188180 1118890 1 0 $X=1188178 $Y=1114950
X790 11258 10299 10952 11331 25 26 MXI2X1 $T=1189100 1089370 1 0 $X=1189098 $Y=1085430
X791 8951 10908 11281 10803 25 26 MXI2X1 $T=1192320 1163170 1 180 $X=1189100 $Y=1162918
X792 11294 11133 10105 11350 25 26 MXI2X1 $T=1190020 1052470 1 0 $X=1190018 $Y=1048530
X793 11331 10299 11143 11284 25 26 MXI2X1 $T=1193240 1089370 1 180 $X=1190020 $Y=1089118
X794 11284 10299 10945 11320 25 26 MXI2X1 $T=1190480 1096750 1 0 $X=1190478 $Y=1092810
X795 11281 140 11388 11021 25 26 MXI2X1 $T=1191400 1163170 1 0 $X=1191398 $Y=1159230
X796 11363 11133 9968 11313 25 26 MXI2X1 $T=1194620 1067230 1 180 $X=1191400 $Y=1066978
X797 11078 11382 11463 11268 25 26 MXI2X1 $T=1196460 1045090 1 0 $X=1196458 $Y=1041150
X798 8951 9196 11499 11196 25 26 MXI2X1 $T=1196460 1133650 1 0 $X=1196458 $Y=1129710
X799 8951 10908 11502 11262 25 26 MXI2X1 $T=1196460 1163170 0 0 $X=1196458 $Y=1162918
X800 11021 140 11414 11173 25 26 MXI2X1 $T=1199680 1163170 0 180 $X=1196460 $Y=1159230
X801 10938 11389 11278 11463 25 26 MXI2X1 $T=1196920 1037710 0 0 $X=1196918 $Y=1037458
X802 11404 11241 11428 11455 25 26 MXI2X1 $T=1196920 1074610 1 0 $X=1196918 $Y=1070670
X803 11439 11030 11265 11351 25 26 MXI2X1 $T=1200140 1067230 0 180 $X=1196920 $Y=1063290
X804 11428 11133 10210 11535 25 26 MXI2X1 $T=1197840 1059850 0 0 $X=1197838 $Y=1059598
X805 8951 11242 11500 11197 25 26 MXI2X1 $T=1197840 1133650 0 0 $X=1197838 $Y=1133398
X806 11261 140 11489 11321 25 26 MXI2X1 $T=1197840 1141030 0 0 $X=1197838 $Y=1140778
X807 11226 140 11501 11198 25 26 MXI2X1 $T=1197840 1155790 0 0 $X=1197838 $Y=1155538
X808 11201 140 11440 11269 25 26 MXI2X1 $T=1201060 1141030 0 180 $X=1197840 $Y=1137090
X809 11467 173 11445 11005 25 26 MXI2X1 $T=1201060 1177930 0 180 $X=1197840 $Y=1173990
X810 11499 140 11574 11201 25 26 MXI2X1 $T=1201980 1133650 1 0 $X=1201978 $Y=1129710
X811 11414 10619 11560 11501 25 26 MXI2X1 $T=1201980 1155790 1 0 $X=1201978 $Y=1151850
X812 11502 140 11594 11373 25 26 MXI2X1 $T=1201980 1163170 0 0 $X=1201978 $Y=1162918
X813 11373 140 11524 11226 25 26 MXI2X1 $T=1205200 1163170 0 180 $X=1201980 $Y=1159230
X814 11268 11382 11506 11629 25 26 MXI2X1 $T=1202900 1045090 1 0 $X=1202898 $Y=1041150
X815 11537 11030 11534 11582 25 26 MXI2X1 $T=1203360 1067230 1 0 $X=1203358 $Y=1063290
X816 11146 173 11585 11467 25 26 MXI2X1 $T=1208880 1170550 0 180 $X=1205660 $Y=1166610
X817 11379 11382 11613 11724 25 26 MXI2X1 $T=1206120 1059850 0 0 $X=1206118 $Y=1059598
X818 10867 140 11733 11261 25 26 MXI2X1 $T=1206120 1133650 0 0 $X=1206118 $Y=1133398
X819 11489 173 11750 11346 25 26 MXI2X1 $T=1206120 1141030 0 0 $X=1206118 $Y=1140778
X820 11388 173 11722 11524 25 26 MXI2X1 $T=1206120 1155790 0 0 $X=1206118 $Y=1155538
X821 11440 173 11589 11489 25 26 MXI2X1 $T=1209340 1141030 0 180 $X=1206120 $Y=1137090
X822 11596 11241 11363 11659 25 26 MXI2X1 $T=1207040 1081990 0 0 $X=1207038 $Y=1081738
X823 11530 173 11727 11669 25 26 MXI2X1 $T=1207500 1126270 0 0 $X=1207498 $Y=1126018
X824 11500 140 11669 10867 25 26 MXI2X1 $T=1207500 1133650 1 0 $X=1207498 $Y=1129710
X825 11501 173 11945 11146 25 26 MXI2X1 $T=1207500 1155790 1 0 $X=1207498 $Y=1151850
X826 11089 173 11643 11594 25 26 MXI2X1 $T=1207500 1163170 0 0 $X=1207498 $Y=1162918
X827 11656 11030 11250 11539 25 26 MXI2X1 $T=1210720 1037710 1 180 $X=1207500 $Y=1037458
X828 11657 11030 11342 11540 25 26 MXI2X1 $T=1210720 1045090 1 180 $X=1207500 $Y=1044838
X829 11658 11030 11330 11439 25 26 MXI2X1 $T=1210720 1067230 1 180 $X=1207500 $Y=1066978
X830 11346 173 11617 11541 25 26 MXI2X1 $T=1210720 1148410 0 180 $X=1207500 $Y=1144470
X831 11524 173 11618 11414 25 26 MXI2X1 $T=1210720 1163170 0 180 $X=1207500 $Y=1159230
X832 11574 173 11861 11733 25 26 MXI2X1 $T=1213020 1133650 1 0 $X=1213018 $Y=1129710
X833 11669 173 11777 11574 25 26 MXI2X1 $T=1213480 1126270 0 0 $X=1213478 $Y=1126018
X834 11594 173 11778 11388 25 26 MXI2X1 $T=1213480 1155790 0 0 $X=1213478 $Y=1155538
X835 11795 11241 11218 11725 25 26 MXI2X1 $T=1216700 1074610 1 180 $X=1213480 $Y=1074358
X836 11796 11389 11608 11739 25 26 MXI2X1 $T=1216700 1081990 0 180 $X=1213480 $Y=1078050
X837 11733 173 11902 11440 25 26 MXI2X1 $T=1213940 1133650 0 0 $X=1213938 $Y=1133398
X838 11658 11389 11398 11796 25 26 MXI2X1 $T=1214860 1074610 1 0 $X=1214858 $Y=1070670
X839 11808 11241 11294 11894 25 26 MXI2X1 $T=1216700 1052470 1 0 $X=1216698 $Y=1048530
X840 11925 11389 11505 11888 25 26 MXI2X1 $T=1222220 1074610 1 180 $X=1219000 $Y=1074358
X841 11956 11241 11686 11912 25 26 MXI2X1 $T=1224060 1074610 0 180 $X=1220840 $Y=1070670
X842 12002 11241 11112 11879 25 26 MXI2X1 $T=1226360 1037710 1 180 $X=1223140 $Y=1037458
X843 11892 11241 11544 11607 25 26 MXI2X1 $T=1225440 1052470 1 0 $X=1225438 $Y=1048530
X844 12040 11241 11965 11565 25 26 MXI2X1 $T=1226360 1030330 0 0 $X=1226358 $Y=1030078
X845 12011 11389 11712 11940 25 26 MXI2X1 $T=1234180 1052470 0 180 $X=1230960 $Y=1048530
X846 11924 11389 11867 12151 25 26 MXI2X1 $T=1232800 1037710 0 0 $X=1232798 $Y=1037458
X847 12063 319 13347 13330 25 26 MXI2X1 $T=1290300 1163170 1 180 $X=1287080 $Y=1162918
X848 12589 319 13641 13632 25 26 MXI2X1 $T=1299960 1141030 0 0 $X=1299958 $Y=1140778
X849 12754 319 13604 13589 25 26 MXI2X1 $T=1299960 1148410 1 0 $X=1299958 $Y=1144470
X850 12754 334 13598 13642 25 26 MXI2X1 $T=1299960 1155790 1 0 $X=1299958 $Y=1151850
X851 12589 335 13643 13633 25 26 MXI2X1 $T=1299960 1155790 0 0 $X=1299958 $Y=1155538
X852 12063 335 13605 13634 25 26 MXI2X1 $T=1299960 1163170 1 0 $X=1299958 $Y=1159230
X853 12258 332 13648 13636 25 26 MXI2X1 $T=1299960 1340290 1 0 $X=1299958 $Y=1336350
X854 13390 319 13594 13638 25 26 MXI2X1 $T=1300420 1273870 0 0 $X=1300418 $Y=1273618
X855 12142 319 13533 13363 25 26 MXI2X1 $T=1304100 1170550 1 180 $X=1300880 $Y=1170298
X856 12050 335 13610 13388 25 26 MXI2X1 $T=1305940 1266490 0 180 $X=1302720 $Y=1262550
X857 13329 319 13682 13584 25 26 MXI2X1 $T=1309160 1273870 1 180 $X=1305940 $Y=1273618
X858 12516 319 13683 13606 25 26 MXI2X1 $T=1309620 1170550 1 180 $X=1306400 $Y=1170298
X859 12024 332 13680 13665 25 26 MXI2X1 $T=1309620 1325530 1 180 $X=1306400 $Y=1325278
X860 230 332 13799 13743 25 26 MXI2X1 $T=1309160 1340290 0 0 $X=1309158 $Y=1340038
X861 12051 343 13674 13658 25 26 MXI2X1 $T=1312840 1288630 1 180 $X=1309620 $Y=1288378
X862 12516 347 13710 13656 25 26 MXI2X1 $T=1313300 1118890 1 180 $X=1310080 $Y=1118638
X863 12516 334 13593 13547 25 26 MXI2X1 $T=1313760 1185310 1 180 $X=1310540 $Y=1185058
X864 13332 319 13713 13650 25 26 MXI2X1 $T=1313760 1244350 1 180 $X=1310540 $Y=1244098
X865 12110 332 13670 13693 25 26 MXI2X1 $T=1313760 1318150 0 180 $X=1310540 $Y=1314210
X866 12792 344 13719 13661 25 26 MXI2X1 $T=1314680 1133650 1 180 $X=1311460 $Y=1133398
X867 12792 319 13657 13583 25 26 MXI2X1 $T=1314680 1170550 1 180 $X=1311460 $Y=1170298
X868 13405 334 13688 13669 25 26 MXI2X1 $T=1311920 1236970 0 0 $X=1311918 $Y=1236718
X869 12589 344 13666 13716 25 26 MXI2X1 $T=1315140 1126270 1 180 $X=1311920 $Y=1126018
X870 12110 343 13664 13747 25 26 MXI2X1 $T=1312380 1303390 1 0 $X=1312378 $Y=1299450
X871 12589 334 13668 13662 25 26 MXI2X1 $T=1312840 1148410 0 0 $X=1312838 $Y=1148158
X872 13390 335 13756 13760 25 26 MXI2X1 $T=1313760 1266490 0 0 $X=1313758 $Y=1266238
X873 12516 350 13812 13840 25 26 MXI2X1 $T=1316980 1118890 1 0 $X=1316978 $Y=1114950
X874 13405 344 13873 13856 25 26 MXI2X1 $T=1316980 1229590 0 0 $X=1316978 $Y=1229338
X875 13332 334 13823 13821 25 26 MXI2X1 $T=1316980 1244350 0 0 $X=1316978 $Y=1244098
X876 12143 334 13777 13781 25 26 MXI2X1 $T=1320200 1192690 0 180 $X=1316980 $Y=1188750
X877 12258 343 13796 351 25 26 MXI2X1 $T=1320200 1340290 0 180 $X=1316980 $Y=1336350
X878 13332 335 13846 13842 25 26 MXI2X1 $T=1317440 1244350 1 0 $X=1317438 $Y=1240410
X879 12063 334 13845 13858 25 26 MXI2X1 $T=1317900 1155790 1 0 $X=1317898 $Y=1151850
X880 12142 334 13787 13841 25 26 MXI2X1 $T=1317900 1163170 0 0 $X=1317898 $Y=1162918
X881 12050 334 13864 13847 25 26 MXI2X1 $T=1317900 1251730 0 0 $X=1317898 $Y=1251478
X882 12050 319 13706 13826 25 26 MXI2X1 $T=1317900 1259110 0 0 $X=1317898 $Y=1258858
X883 12024 353 13798 13850 25 26 MXI2X1 $T=1317900 1332910 1 0 $X=1317898 $Y=1328970
X884 12516 344 13773 13801 25 26 MXI2X1 $T=1321120 1133650 0 180 $X=1317900 $Y=1129710
X885 12754 335 13809 13774 25 26 MXI2X1 $T=1321120 1148410 1 180 $X=1317900 $Y=1148158
X886 13390 334 13772 13771 25 26 MXI2X1 $T=1321120 1273870 0 180 $X=1317900 $Y=1269930
X887 13329 335 13778 13733 25 26 MXI2X1 $T=1321120 1281250 0 180 $X=1317900 $Y=1277310
X888 12024 343 13776 13794 25 26 MXI2X1 $T=1321120 1325530 0 180 $X=1317900 $Y=1321590
X889 12792 350 13820 13805 25 26 MXI2X1 $T=1318360 1104130 0 0 $X=1318358 $Y=1103878
X890 12143 319 13759 13872 25 26 MXI2X1 $T=1318360 1222210 1 0 $X=1318358 $Y=1218270
X891 230 353 13789 13874 25 26 MXI2X1 $T=1318360 1347670 1 0 $X=1318358 $Y=1343730
X892 12143 335 13795 13822 25 26 MXI2X1 $T=1318820 1200070 0 0 $X=1318818 $Y=1199818
X893 12516 335 13817 13815 25 26 MXI2X1 $T=1322500 1185310 1 180 $X=1319280 $Y=1185058
X894 12039 319 13818 13752 25 26 MXI2X1 $T=1322500 1214830 0 180 $X=1319280 $Y=1210890
X895 13405 350 13829 13686 25 26 MXI2X1 $T=1322960 1236970 0 180 $X=1319740 $Y=1233030
X896 12110 353 13827 13762 25 26 MXI2X1 $T=1322960 1318150 0 180 $X=1319740 $Y=1314210
X897 12110 358 13861 13878 25 26 MXI2X1 $T=1320660 1310770 0 0 $X=1320658 $Y=1310518
X898 12143 347 13969 13770 25 26 MXI2X1 $T=1321580 1192690 1 0 $X=1321578 $Y=1188750
X899 13329 334 13848 356 25 26 MXI2X1 $T=1324800 1288630 1 180 $X=1321580 $Y=1288378
X900 13390 344 13917 13921 25 26 MXI2X1 $T=1323880 1251730 0 0 $X=1323878 $Y=1251478
X901 12754 344 13802 13855 25 26 MXI2X1 $T=1327100 1133650 1 180 $X=1323880 $Y=1133398
X902 12258 353 13862 13922 25 26 MXI2X1 $T=1324800 1347670 1 0 $X=1324798 $Y=1343730
X903 13390 347 13898 13910 25 26 MXI2X1 $T=1326640 1259110 0 0 $X=1326638 $Y=1258858
X904 12051 353 13909 13849 25 26 MXI2X1 $T=1326640 1310770 1 0 $X=1326638 $Y=1306830
X905 12792 334 13825 13908 25 26 MXI2X1 $T=1328020 1185310 0 0 $X=1328018 $Y=1185058
X906 12039 334 13830 13814 25 26 MXI2X1 $T=1328020 1214830 1 0 $X=1328018 $Y=1210890
X907 13405 347 13899 13959 25 26 MXI2X1 $T=1328940 1222210 1 0 $X=1328938 $Y=1218270
X908 12142 335 13987 14003 25 26 MXI2X1 $T=1330780 1177930 1 0 $X=1330778 $Y=1173990
X909 13405 382 14112 13970 25 26 MXI2X1 $T=1332620 1236970 0 0 $X=1332618 $Y=1236718
X910 12051 384 13979 14002 25 26 MXI2X1 $T=1333540 1296010 0 0 $X=1333538 $Y=1295758
X911 12516 382 13950 13857 25 26 MXI2X1 $T=1336760 1126270 0 180 $X=1333540 $Y=1122330
X912 12589 382 13994 14024 25 26 MXI2X1 $T=1334460 1111510 1 0 $X=1334458 $Y=1107570
X913 12142 344 14026 14027 25 26 MXI2X1 $T=1334460 1133650 1 0 $X=1334458 $Y=1129710
X914 12143 382 14030 14029 25 26 MXI2X1 $T=1334460 1185310 0 0 $X=1334458 $Y=1185058
X915 13332 347 13999 13806 25 26 MXI2X1 $T=1334460 1222210 1 0 $X=1334458 $Y=1218270
X916 12024 384 14013 14020 25 26 MXI2X1 $T=1334460 1325530 0 0 $X=1334458 $Y=1325278
X917 12754 382 13854 13751 25 26 MXI2X1 $T=1337680 1111510 1 180 $X=1334460 $Y=1111258
X918 12110 391 13980 13946 25 26 MXI2X1 $T=1337680 1303390 1 180 $X=1334460 $Y=1303138
X919 12039 350 14043 14016 25 26 MXI2X1 $T=1334920 1200070 0 0 $X=1334918 $Y=1199818
X920 12589 350 14010 13967 25 26 MXI2X1 $T=1335380 1148410 0 0 $X=1335378 $Y=1148158
X921 12143 344 14051 14028 25 26 MXI2X1 $T=1335380 1185310 1 0 $X=1335378 $Y=1181370
X922 12039 344 14044 14064 25 26 MXI2X1 $T=1335380 1214830 1 0 $X=1335378 $Y=1210890
X923 13329 347 14012 14034 25 26 MXI2X1 $T=1335380 1273870 1 0 $X=1335378 $Y=1269930
X924 12589 347 13863 13766 25 26 MXI2X1 $T=1338600 1133650 1 180 $X=1335380 $Y=1133398
X925 12063 344 13996 13758 25 26 MXI2X1 $T=1338600 1170550 1 180 $X=1335380 $Y=1170298
X926 13329 350 13978 13930 25 26 MXI2X1 $T=1338600 1281250 0 180 $X=1335380 $Y=1277310
X927 13390 350 14089 14068 25 26 MXI2X1 $T=1335840 1266490 0 0 $X=1335838 $Y=1266238
X928 12754 350 13941 14062 25 26 MXI2X1 $T=1336760 1104130 0 0 $X=1336758 $Y=1103878
X929 12039 335 13956 14088 25 26 MXI2X1 $T=1336760 1207450 1 0 $X=1336758 $Y=1203510
X930 12051 393 14059 14090 25 26 MXI2X1 $T=1336760 1296010 0 0 $X=1336758 $Y=1295758
X931 12024 358 14056 14045 25 26 MXI2X1 $T=1336760 1325530 1 0 $X=1336758 $Y=1321590
X932 12258 384 13990 14006 25 26 MXI2X1 $T=1340900 1332910 1 180 $X=1337680 $Y=1332658
X933 13390 382 14049 14052 25 26 MXI2X1 $T=1343200 1251730 1 180 $X=1339980 $Y=1251478
X934 12063 350 13982 13951 25 26 MXI2X1 $T=1340440 1155790 1 0 $X=1340438 $Y=1151850
X935 12258 393 14106 14104 25 26 MXI2X1 $T=1340900 1332910 0 0 $X=1340898 $Y=1332658
X936 13329 344 14014 14005 25 26 MXI2X1 $T=1344120 1281250 0 180 $X=1340900 $Y=1277310
X937 12024 391 14050 13900 25 26 MXI2X1 $T=1344120 1310770 1 180 $X=1340900 $Y=1310518
X938 12050 347 14117 14122 25 26 MXI2X1 $T=1343200 1251730 0 0 $X=1343198 $Y=1251478
X939 12792 382 14115 13813 25 26 MXI2X1 $T=1348260 1104130 1 180 $X=1345040 $Y=1103878
X940 12039 347 14084 13952 25 26 MXI2X1 $T=1348260 1207450 0 180 $X=1345040 $Y=1203510
X941 12024 393 14118 14046 25 26 MXI2X1 $T=1348260 1325530 0 180 $X=1345040 $Y=1321590
X942 12051 358 14036 14129 25 26 MXI2X1 $T=1346420 1310770 0 0 $X=1346418 $Y=1310518
X943 13329 382 14105 14004 25 26 MXI2X1 $T=1349640 1281250 0 180 $X=1346420 $Y=1277310
X944 14131 315 13114 14175 25 26 MXI2X1 $T=1347340 1244350 1 0 $X=1347338 $Y=1240410
X945 13332 344 14113 13867 25 26 MXI2X1 $T=1350560 1229590 1 180 $X=1347340 $Y=1229338
X946 12050 382 14134 14092 25 26 MXI2X1 $T=1351480 1251730 0 180 $X=1348260 $Y=1247790
X947 12063 347 13955 14094 25 26 MXI2X1 $T=1351940 1163170 0 180 $X=1348720 $Y=1159230
X948 12051 391 14066 14100 25 26 MXI2X1 $T=1352860 1288630 1 180 $X=1349640 $Y=1288378
X949 14174 53 12758 14207 25 26 MXI2X1 $T=1351480 1185310 1 0 $X=1351478 $Y=1181370
X950 14140 53 12369 14217 25 26 MXI2X1 $T=1352400 1177930 0 0 $X=1352398 $Y=1177678
X951 14192 83 12146 14218 25 26 MXI2X1 $T=1352400 1185310 0 0 $X=1352398 $Y=1185058
X952 14194 83 12946 14221 25 26 MXI2X1 $T=1352400 1281250 0 0 $X=1352398 $Y=1280998
X953 13332 382 14193 14085 25 26 MXI2X1 $T=1355620 1229590 0 180 $X=1352400 $Y=1225650
X954 12063 382 14167 14234 25 26 MXI2X1 $T=1353780 1177930 1 0 $X=1353778 $Y=1173990
X955 12142 382 14185 14095 25 26 MXI2X1 $T=1357000 1111510 0 180 $X=1353780 $Y=1107570
X956 14211 83 12651 14236 25 26 MXI2X1 $T=1354240 1236970 0 0 $X=1354238 $Y=1236718
X957 12792 411 14209 14155 25 26 MXI2X1 $T=1357460 1170550 0 180 $X=1354240 $Y=1166610
X958 12754 347 14054 14148 25 26 MXI2X1 $T=1354700 1133650 0 0 $X=1354698 $Y=1133398
X959 407 425 12165 404 25 26 MXI2X1 $T=1357920 1347670 1 180 $X=1354700 $Y=1347418
X960 12110 393 14170 14213 25 26 MXI2X1 $T=1358840 1296010 1 180 $X=1355620 $Y=1295758
X961 12589 409 14189 14269 25 26 MXI2X1 $T=1356080 1111510 0 0 $X=1356078 $Y=1111258
X962 12792 409 14368 14183 25 26 MXI2X1 $T=1356080 1126270 1 0 $X=1356078 $Y=1122330
X963 12039 382 14263 14041 25 26 MXI2X1 $T=1356080 1200070 0 0 $X=1356078 $Y=1199818
X964 14241 408 11468 14265 25 26 MXI2X1 $T=1357000 1340290 0 0 $X=1356998 $Y=1340038
X965 12143 350 14238 14297 25 26 MXI2X1 $T=1358380 1185310 0 0 $X=1358378 $Y=1185058
X966 14232 425 11528 14322 25 26 MXI2X1 $T=1361600 1207450 1 0 $X=1361598 $Y=1203510
X967 12050 344 14311 14204 25 26 MXI2X1 $T=1362060 1259110 0 0 $X=1362058 $Y=1258858
X968 12516 409 14223 14336 25 26 MXI2X1 $T=1362520 1133650 0 0 $X=1362518 $Y=1133398
X969 14248 53 12501 14342 25 26 MXI2X1 $T=1362520 1177930 1 0 $X=1362518 $Y=1173990
X970 14305 83 12864 14348 25 26 MXI2X1 $T=1362520 1273870 0 0 $X=1362518 $Y=1273618
X971 14308 408 11214 14361 25 26 MXI2X1 $T=1362520 1325530 0 0 $X=1362518 $Y=1325278
X972 12589 427 14304 14188 25 26 MXI2X1 $T=1365740 1111510 0 180 $X=1362520 $Y=1107570
X973 14321 408 12255 14352 25 26 MXI2X1 $T=1363900 1185310 0 0 $X=1363898 $Y=1185058
X974 14350 408 11516 14272 25 26 MXI2X1 $T=1367120 1303390 1 180 $X=1363900 $Y=1303138
X975 12050 350 14334 14130 25 26 MXI2X1 $T=1367580 1244350 1 180 $X=1364360 $Y=1244098
X976 12142 350 14300 14323 25 26 MXI2X1 $T=1364820 1118890 1 0 $X=1364818 $Y=1114950
X977 12039 433 14343 14327 25 26 MXI2X1 $T=1368040 1200070 1 180 $X=1364820 $Y=1199818
X978 14356 408 13188 14329 25 26 MXI2X1 $T=1368040 1229590 1 180 $X=1364820 $Y=1229338
X979 12039 409 14370 14267 25 26 MXI2X1 $T=1365740 1214830 1 0 $X=1365738 $Y=1210890
X980 12051 436 14222 14338 25 26 MXI2X1 $T=1369420 1310770 1 180 $X=1366200 $Y=1310518
X981 14383 408 11296 14359 25 26 MXI2X1 $T=1370340 1318150 0 180 $X=1367120 $Y=1314210
X982 12589 433 14395 14399 25 26 MXI2X1 $T=1368040 1141030 1 0 $X=1368038 $Y=1137090
X983 13405 427 14384 14344 25 26 MXI2X1 $T=1368040 1244350 0 0 $X=1368038 $Y=1244098
X984 14366 425 12359 14402 25 26 MXI2X1 $T=1368040 1296010 1 0 $X=1368038 $Y=1292070
X985 14251 53 12922 14417 25 26 MXI2X1 $T=1368500 1259110 0 0 $X=1368498 $Y=1258858
X986 12754 427 14419 14425 25 26 MXI2X1 $T=1368960 1104130 0 0 $X=1368958 $Y=1103878
X987 12792 427 14426 14420 25 26 MXI2X1 $T=1368960 1111510 1 0 $X=1368958 $Y=1107570
X988 12143 411 14396 14428 25 26 MXI2X1 $T=1368960 1185310 1 0 $X=1368958 $Y=1181370
X989 12039 411 14429 14422 25 26 MXI2X1 $T=1368960 1200070 1 0 $X=1368958 $Y=1196130
X990 14382 83 12921 14430 25 26 MXI2X1 $T=1368960 1222210 1 0 $X=1368958 $Y=1218270
X991 14371 425 12156 14431 25 26 MXI2X1 $T=1368960 1325530 0 0 $X=1368958 $Y=1325278
X992 14386 408 11646 14441 25 26 MXI2X1 $T=1369420 1214830 0 0 $X=1369418 $Y=1214578
X993 14392 83 12014 14468 25 26 MXI2X1 $T=1369880 1177930 1 0 $X=1369878 $Y=1173990
X994 12110 436 14469 14314 25 26 MXI2X1 $T=1369880 1281250 1 0 $X=1369878 $Y=1277310
X995 14390 425 11661 14450 25 26 MXI2X1 $T=1369880 1310770 1 0 $X=1369878 $Y=1306830
X996 14379 425 12164 14471 25 26 MXI2X1 $T=1369880 1318150 0 0 $X=1369878 $Y=1317898
X997 12024 436 14460 14442 25 26 MXI2X1 $T=1369880 1325530 1 0 $X=1369878 $Y=1321590
X998 12754 411 14447 14452 25 26 MXI2X1 $T=1371260 1141030 1 0 $X=1371258 $Y=1137090
X999 13390 411 14473 14345 25 26 MXI2X1 $T=1371260 1266490 0 0 $X=1371258 $Y=1266238
X1000 12516 427 14421 14374 25 26 MXI2X1 $T=1374480 1126270 0 180 $X=1371260 $Y=1122330
X1001 12051 437 14470 14378 25 26 MXI2X1 $T=1373100 1303390 0 0 $X=1373098 $Y=1303138
X1002 12143 433 14443 14381 25 26 MXI2X1 $T=1376320 1185310 0 180 $X=1373100 $Y=1181370
X1003 13390 409 14459 14364 25 26 MXI2X1 $T=1376780 1251730 0 180 $X=1373560 $Y=1247790
X1004 12754 409 14462 14514 25 26 MXI2X1 $T=1375400 1111510 0 0 $X=1375398 $Y=1111258
X1005 14478 83 12368 14515 25 26 MXI2X1 $T=1375400 1177930 1 0 $X=1375398 $Y=1173990
X1006 12258 436 14363 14461 25 26 MXI2X1 $T=1375400 1340290 0 0 $X=1375398 $Y=1340038
X1007 12516 433 14511 14398 25 26 MXI2X1 $T=1382760 1126270 0 180 $X=1379540 $Y=1122330
X1008 13329 411 14512 14477 25 26 MXI2X1 $T=1382760 1266490 1 180 $X=1379540 $Y=1266238
X1009 12024 437 14423 14451 25 26 MXI2X1 $T=1382760 1310770 1 180 $X=1379540 $Y=1310518
X1010 14520 425 11443 14559 25 26 MXI2X1 $T=1380460 1170550 0 0 $X=1380458 $Y=1170298
X1011 14388 430 11558 14594 25 26 MXI2X1 $T=1380460 1288630 0 0 $X=1380458 $Y=1288378
X1012 12142 411 14492 14508 25 26 MXI2X1 $T=1383680 1155790 0 180 $X=1380460 $Y=1151850
X1013 14516 430 12392 14565 25 26 MXI2X1 $T=1380920 1192690 0 0 $X=1380918 $Y=1192438
X1014 14517 430 11581 14554 25 26 MXI2X1 $T=1380920 1251730 0 0 $X=1380918 $Y=1251478
X1015 12754 433 14522 14456 25 26 MXI2X1 $T=1384140 1111510 1 180 $X=1380920 $Y=1111258
X1016 12258 437 14504 14349 25 26 MXI2X1 $T=1384140 1332910 0 180 $X=1380920 $Y=1328970
X1017 13405 409 14545 14444 25 26 MXI2X1 $T=1381380 1214830 0 0 $X=1381378 $Y=1214578
X1018 13405 411 14362 14249 25 26 MXI2X1 $T=1384600 1236970 0 180 $X=1381380 $Y=1233030
X1019 14521 425 11673 14560 25 26 MXI2X1 $T=1381840 1259110 0 0 $X=1381838 $Y=1258858
X1020 12516 411 14506 14303 25 26 MXI2X1 $T=1385060 1155790 1 180 $X=1381840 $Y=1155538
X1021 12143 427 14538 14448 25 26 MXI2X1 $T=1385060 1177930 1 180 $X=1381840 $Y=1177678
X1022 13390 427 14541 14486 25 26 MXI2X1 $T=1385060 1259110 0 180 $X=1381840 $Y=1255170
X1023 12110 448 14481 14562 25 26 MXI2X1 $T=1384140 1296010 0 0 $X=1384138 $Y=1295758
X1024 14566 425 11622 14598 25 26 MXI2X1 $T=1385520 1170550 0 0 $X=1385518 $Y=1170298
X1025 12143 409 14584 14615 25 26 MXI2X1 $T=1385980 1200070 1 0 $X=1385978 $Y=1196130
X1026 14570 425 11800 14616 25 26 MXI2X1 $T=1385980 1214830 0 0 $X=1385978 $Y=1214578
X1027 12050 411 14585 14472 25 26 MXI2X1 $T=1385980 1244350 1 0 $X=1385978 $Y=1240410
X1028 13329 409 14588 14572 25 26 MXI2X1 $T=1385980 1266490 0 0 $X=1385978 $Y=1266238
X1029 12051 447 14601 14608 25 26 MXI2X1 $T=1385980 1310770 1 0 $X=1385978 $Y=1306830
X1030 12792 433 14551 14457 25 26 MXI2X1 $T=1389200 1133650 1 180 $X=1385980 $Y=1133398
X1031 12589 411 14377 14266 25 26 MXI2X1 $T=1389200 1141030 1 180 $X=1385980 $Y=1140778
X1032 13329 427 14577 14549 25 26 MXI2X1 $T=1389200 1281250 0 180 $X=1385980 $Y=1277310
X1033 13332 411 14576 14488 25 26 MXI2X1 $T=1389660 1236970 0 180 $X=1386440 $Y=1233030
X1034 12050 409 14606 14617 25 26 MXI2X1 $T=1386900 1251730 0 0 $X=1386898 $Y=1251478
X1035 12024 448 14659 14621 25 26 MXI2X1 $T=1386900 1318150 0 0 $X=1386898 $Y=1317898
X1036 230 448 14602 14613 25 26 MXI2X1 $T=1386900 1347670 1 0 $X=1386898 $Y=1343730
X1037 13332 409 14568 14482 25 26 MXI2X1 $T=1390120 1222210 1 180 $X=1386900 $Y=1221958
X1038 12063 427 14583 14685 25 26 MXI2X1 $T=1388280 1104130 0 0 $X=1388278 $Y=1103878
X1039 12039 453 14605 14696 25 26 MXI2X1 $T=1388280 1214830 1 0 $X=1388278 $Y=1210890
X1040 12142 433 14603 14573 25 26 MXI2X1 $T=1391500 1118890 0 180 $X=1388280 $Y=1114950
X1041 230 450 14641 14660 25 26 MXI2X1 $T=1388740 1340290 0 0 $X=1388738 $Y=1340038
X1042 12063 14639 14609 14574 25 26 MXI2X1 $T=1391960 1170550 1 180 $X=1388740 $Y=1170298
X1043 12024 452 14631 14646 25 26 MXI2X1 $T=1389200 1310770 1 0 $X=1389198 $Y=1306830
X1044 12143 14639 14627 14612 25 26 MXI2X1 $T=1392880 1185310 1 180 $X=1389660 $Y=1185058
X1045 13329 433 14667 14624 25 26 MXI2X1 $T=1390120 1266490 0 0 $X=1390118 $Y=1266238
X1046 12051 452 14618 14676 25 26 MXI2X1 $T=1390120 1296010 1 0 $X=1390118 $Y=1292070
X1047 13390 433 14630 14569 25 26 MXI2X1 $T=1393340 1266490 0 180 $X=1390120 $Y=1262550
X1048 12110 452 14665 14620 25 26 MXI2X1 $T=1390580 1310770 0 0 $X=1390578 $Y=1310518
X1049 13329 453 14712 14713 25 26 MXI2X1 $T=1391500 1281250 1 0 $X=1391498 $Y=1277310
X1050 12110 447 14625 14519 25 26 MXI2X1 $T=1395180 1288630 0 180 $X=1391960 $Y=1284690
X1051 13332 427 14670 14548 25 26 MXI2X1 $T=1396100 1222210 1 180 $X=1392880 $Y=1221958
X1052 12039 14639 14645 14592 25 26 MXI2X1 $T=1397940 1200070 1 180 $X=1394720 $Y=1199818
X1053 12063 411 14729 14633 25 26 MXI2X1 $T=1396100 1141030 1 0 $X=1396098 $Y=1137090
X1054 12051 448 14747 14668 25 26 MXI2X1 $T=1397020 1303390 0 0 $X=1397018 $Y=1303138
X1055 12142 427 14694 14537 25 26 MXI2X1 $T=1400240 1104130 1 180 $X=1397020 $Y=1103878
X1056 12063 433 14695 14600 25 26 MXI2X1 $T=1400240 1118890 0 180 $X=1397020 $Y=1114950
X1057 12142 14639 14587 14397 25 26 MXI2X1 $T=1400240 1185310 0 180 $X=1397020 $Y=1181370
X1058 12050 427 14509 14610 25 26 MXI2X1 $T=1400240 1244350 1 180 $X=1397020 $Y=1244098
X1059 12142 453 14557 14487 25 26 MXI2X1 $T=1401160 1148410 1 180 $X=1397940 $Y=1148158
X1060 13332 433 14703 14593 25 26 MXI2X1 $T=1401620 1222210 1 180 $X=1398400 $Y=1221958
X1061 12039 427 14701 14575 25 26 MXI2X1 $T=1399320 1192690 0 0 $X=1399318 $Y=1192438
X1062 12024 447 14679 14582 25 26 MXI2X1 $T=1399320 1325530 0 0 $X=1399318 $Y=1325278
X1063 12258 448 14680 14578 25 26 MXI2X1 $T=1399320 1332910 1 0 $X=1399318 $Y=1328970
X1064 12792 14639 14708 14682 25 26 MXI2X1 $T=1402540 1177930 0 180 $X=1399320 $Y=1173990
X1065 13405 433 14711 14635 25 26 MXI2X1 $T=1402540 1236970 1 180 $X=1399320 $Y=1236718
X1066 12063 14773 14738 14643 25 26 MXI2X1 $T=1405760 1155790 1 180 $X=1402540 $Y=1155538
X1067 12754 453 14767 14734 25 26 MXI2X1 $T=1403460 1133650 0 0 $X=1403458 $Y=1133398
X1068 12516 14639 14769 14781 25 26 MXI2X1 $T=1403460 1185310 1 0 $X=1403458 $Y=1181370
X1069 13390 453 14746 14739 25 26 MXI2X1 $T=1406680 1266490 0 180 $X=1403460 $Y=1262550
X1070 12050 453 14684 14778 25 26 MXI2X1 $T=1404380 1281250 0 0 $X=1404378 $Y=1280998
X1071 13332 14773 14640 14706 25 26 MXI2X1 $T=1407600 1222210 0 180 $X=1404380 $Y=1218270
X1072 13405 453 14771 14697 25 26 MXI2X1 $T=1407600 1244350 1 180 $X=1404380 $Y=1244098
X1073 12050 14639 14765 14733 25 26 MXI2X1 $T=1407600 1259110 0 180 $X=1404380 $Y=1255170
X1074 12142 409 14779 14761 25 26 MXI2X1 $T=1408980 1118890 0 180 $X=1405760 $Y=1114950
X1075 12063 409 14748 14662 25 26 MXI2X1 $T=1408980 1126270 1 180 $X=1405760 $Y=1126018
X1076 12142 14773 14730 14637 25 26 MXI2X1 $T=1408980 1141030 0 180 $X=1405760 $Y=1137090
X1077 12792 14773 14772 14675 25 26 MXI2X1 $T=1408980 1148410 1 180 $X=1405760 $Y=1148158
X1078 12258 452 14666 14683 25 26 MXI2X1 $T=1408980 1332910 1 180 $X=1405760 $Y=1332658
X1079 12143 453 14709 14809 25 26 MXI2X1 $T=1406220 1207450 1 0 $X=1406218 $Y=1203510
X1080 12516 14773 14832 14796 25 26 MXI2X1 $T=1409440 1177930 0 0 $X=1409438 $Y=1177678
X1081 12051 470 14808 14886 25 26 MXI2X1 $T=1409900 1288630 0 0 $X=1409898 $Y=1288378
X1082 13405 14773 14815 14777 25 26 MXI2X1 $T=1413120 1244350 1 180 $X=1409900 $Y=1244098
X1083 13332 453 14836 14817 25 26 MXI2X1 $T=1414040 1222210 0 180 $X=1410820 $Y=1218270
X1084 12063 453 14841 14786 25 26 MXI2X1 $T=1415420 1163170 1 180 $X=1412200 $Y=1162918
X1085 14867 473 14859 14766 25 26 MXI2X1 $T=1417260 1118890 0 180 $X=1414040 $Y=1114950
X1086 12792 453 14854 14768 25 26 MXI2X1 $T=1417260 1148410 1 180 $X=1414040 $Y=1148158
X1087 12110 470 14775 14853 25 26 MXI2X1 $T=1417260 1310770 1 180 $X=1414040 $Y=1310518
X1088 12258 470 14861 14782 25 26 MXI2X1 $T=1417260 1332910 1 180 $X=1414040 $Y=1332658
X1089 12516 453 14888 14806 25 26 MXI2X1 $T=1415420 1177930 1 0 $X=1415418 $Y=1173990
X1090 13332 14639 14873 14849 25 26 MXI2X1 $T=1415420 1229590 1 0 $X=1415418 $Y=1225650
X1091 13390 14639 14850 14920 25 26 MXI2X1 $T=1415420 1244350 0 0 $X=1415418 $Y=1244098
X1092 12050 450 14882 14802 25 26 MXI2X1 $T=1415420 1273870 1 0 $X=1415418 $Y=1269930
X1093 12110 450 14895 14835 25 26 MXI2X1 $T=1415420 1303390 1 0 $X=1415418 $Y=1299450
X1094 12143 14773 14856 14770 25 26 MXI2X1 $T=1418640 1192690 1 180 $X=1415420 $Y=1192438
X1095 12039 14773 14866 14844 25 26 MXI2X1 $T=1418640 1207450 0 180 $X=1415420 $Y=1203510
X1096 14879 473 14852 14755 25 26 MXI2X1 $T=1418640 1214830 0 180 $X=1415420 $Y=1210890
X1097 12024 470 14846 14754 25 26 MXI2X1 $T=1418640 1325530 0 180 $X=1415420 $Y=1321590
X1098 12754 14773 14855 14762 25 26 MXI2X1 $T=1419560 1133650 0 180 $X=1416340 $Y=1129710
X1099 12039 475 14759 14634 25 26 MXI2X1 $T=1420020 1222210 0 180 $X=1416800 $Y=1218270
X1100 14917 14921 14891 14864 25 26 MXI2X1 $T=1422320 1259110 0 180 $X=1419100 $Y=1255170
X1101 12589 453 14799 14735 25 26 MXI2X1 $T=1420020 1141030 1 0 $X=1420018 $Y=1137090
X1102 12050 480 14880 14792 25 26 MXI2X1 $T=1423240 1273870 1 180 $X=1420020 $Y=1273618
X1103 14929 474 14900 476 25 26 MXI2X1 $T=1423700 1347670 0 180 $X=1420480 $Y=1343730
X1104 13405 14639 14916 14862 25 26 MXI2X1 $T=1424160 1236970 1 180 $X=1420940 $Y=1236718
X1105 14937 480 14899 14834 25 26 MXI2X1 $T=1425080 1288630 1 180 $X=1421860 $Y=1288378
X1106 14926 473 14912 14636 25 26 MXI2X1 $T=1425080 1303390 0 180 $X=1421860 $Y=1299450
X1107 14926 14773 14863 14760 25 26 MXI2X1 $T=1425080 1318150 1 180 $X=1421860 $Y=1317898
X1108 12142 475 14956 14994 25 26 MXI2X1 $T=1422780 1177930 1 0 $X=1422778 $Y=1173990
X1109 12063 475 14963 14954 25 26 MXI2X1 $T=1422780 1185310 0 0 $X=1422778 $Y=1185058
X1110 13329 14773 14970 14881 25 26 MXI2X1 $T=1422780 1288630 1 0 $X=1422778 $Y=1284690
X1111 14867 14936 14925 14928 25 26 MXI2X1 $T=1426000 1155790 0 180 $X=1422780 $Y=1151850
X1112 12589 14639 14877 14795 25 26 MXI2X1 $T=1426000 1163170 0 180 $X=1422780 $Y=1159230
X1113 14879 14921 14964 15013 25 26 MXI2X1 $T=1423240 1222210 0 0 $X=1423238 $Y=1221958
X1114 13390 14773 14947 14885 25 26 MXI2X1 $T=1423240 1266490 0 0 $X=1423238 $Y=1266238
X1115 12051 481 14948 15031 25 26 MXI2X1 $T=1423240 1296010 0 0 $X=1423238 $Y=1295758
X1116 14955 473 14892 14816 25 26 MXI2X1 $T=1426460 1192690 1 180 $X=1423240 $Y=1192438
X1117 12110 480 14932 14851 25 26 MXI2X1 $T=1426460 1318150 0 180 $X=1423240 $Y=1314210
X1118 14966 473 14943 14858 25 26 MXI2X1 $T=1427380 1118890 1 180 $X=1424160 $Y=1118638
X1119 14955 14921 14951 14889 25 26 MXI2X1 $T=1427840 1200070 1 180 $X=1424620 $Y=1199818
X1120 14955 14936 14915 14939 25 26 MXI2X1 $T=1427840 1207450 1 180 $X=1424620 $Y=1207198
X1121 12589 14773 14927 15012 25 26 MXI2X1 $T=1426460 1141030 1 0 $X=1426458 $Y=1137090
X1122 13405 473 14972 14930 25 26 MXI2X1 $T=1430140 1236970 1 180 $X=1426920 $Y=1236718
X1123 230 481 14983 14969 25 26 MXI2X1 $T=1427380 1347670 0 0 $X=1427378 $Y=1347418
X1124 12110 481 14984 14945 25 26 MXI2X1 $T=1431520 1303390 0 180 $X=1428300 $Y=1299450
X1125 12024 481 14982 14938 25 26 MXI2X1 $T=1431520 1318150 1 180 $X=1428300 $Y=1317898
X1126 14992 473 14986 14944 25 26 MXI2X1 $T=1431980 1133650 1 180 $X=1428760 $Y=1133398
X1127 13332 473 14991 14923 25 26 MXI2X1 $T=1433360 1229590 1 180 $X=1430140 $Y=1229338
X1128 12050 475 14933 15019 25 26 MXI2X1 $T=1430600 1251730 1 0 $X=1430598 $Y=1247790
X1129 12024 489 14965 15027 25 26 MXI2X1 $T=1431060 1332910 1 0 $X=1431058 $Y=1328970
X1130 14937 489 14996 14952 25 26 MXI2X1 $T=1434280 1288630 0 180 $X=1431060 $Y=1284690
X1131 14929 473 14997 14941 25 26 MXI2X1 $T=1434280 1340290 0 180 $X=1431060 $Y=1336350
X1132 12792 475 14931 14957 25 26 MXI2X1 $T=1431520 1185310 0 0 $X=1431518 $Y=1185058
X1133 14913 14921 14980 14976 25 26 MXI2X1 $T=1434740 1155790 0 180 $X=1431520 $Y=1151850
X1134 14867 14921 14878 14950 25 26 MXI2X1 $T=1434740 1163170 0 180 $X=1431520 $Y=1159230
X1135 15020 473 14990 14914 25 26 MXI2X1 $T=1434740 1177930 0 180 $X=1431520 $Y=1173990
X1136 12143 475 14987 14981 25 26 MXI2X1 $T=1432440 1214830 1 0 $X=1432438 $Y=1210890
X1137 15022 493 14960 15014 25 26 MXI2X1 $T=1435660 1310770 0 180 $X=1432440 $Y=1306830
X1138 14913 14936 14979 14922 25 26 MXI2X1 $T=1436120 1141030 0 180 $X=1432900 $Y=1137090
X1139 13329 473 14973 15040 25 26 MXI2X1 $T=1433820 1281250 1 0 $X=1433818 $Y=1277310
X1140 14993 473 15024 14949 25 26 MXI2X1 $T=1437040 1118890 0 180 $X=1433820 $Y=1114950
X1141 14926 493 15044 15023 25 26 MXI2X1 $T=1434740 1318150 0 0 $X=1434738 $Y=1317898
X1142 12258 481 14971 15041 25 26 MXI2X1 $T=1436120 1340290 1 0 $X=1436118 $Y=1336350
X1143 15053 473 15026 14946 25 26 MXI2X1 $T=1439340 1259110 0 180 $X=1436120 $Y=1255170
X1144 14917 14936 15052 15032 25 26 MXI2X1 $T=1436580 1244350 1 0 $X=1436578 $Y=1240410
X1145 14879 14936 15042 14958 25 26 MXI2X1 $T=1439800 1229590 0 180 $X=1436580 $Y=1225650
X1146 14955 15057 15116 15129 25 26 MXI2X1 $T=1437500 1185310 0 0 $X=1437498 $Y=1185058
X1147 14937 493 15087 15081 25 26 MXI2X1 $T=1437960 1303390 1 0 $X=1437958 $Y=1299450
X1148 14867 15057 14968 15030 25 26 MXI2X1 $T=1441180 1118890 1 180 $X=1437960 $Y=1118638
X1149 14937 496 15060 15086 25 26 MXI2X1 $T=1438420 1273870 0 0 $X=1438418 $Y=1273618
X1150 14913 15057 15122 14962 25 26 MXI2X1 $T=1438880 1126270 0 0 $X=1438878 $Y=1126018
X1151 12516 475 14967 15034 25 26 MXI2X1 $T=1438880 1177930 1 0 $X=1438878 $Y=1173990
X1152 14867 15075 15055 14919 25 26 MXI2X1 $T=1442100 1163170 0 180 $X=1438880 $Y=1159230
X1153 14955 15075 15064 15056 25 26 MXI2X1 $T=1442100 1200070 0 180 $X=1438880 $Y=1196130
X1154 497 489 15074 14977 25 26 MXI2X1 $T=1442560 1347670 0 180 $X=1439340 $Y=1343730
X1155 14913 15075 15165 15080 25 26 MXI2X1 $T=1440260 1141030 0 0 $X=1440258 $Y=1140778
X1156 12754 475 15091 15058 25 26 MXI2X1 $T=1440260 1185310 1 0 $X=1440258 $Y=1181370
X1157 14879 15075 15092 15120 25 26 MXI2X1 $T=1440260 1207450 0 0 $X=1440258 $Y=1207198
X1158 14929 493 15050 15125 25 26 MXI2X1 $T=1440720 1325530 0 0 $X=1440718 $Y=1325278
X1159 14955 15131 15084 15083 25 26 MXI2X1 $T=1444400 1229590 0 180 $X=1441180 $Y=1225650
X1160 15022 489 15124 14953 25 26 MXI2X1 $T=1441640 1318150 0 0 $X=1441638 $Y=1317898
X1161 14879 15057 15146 15123 25 26 MXI2X1 $T=1444400 1229590 1 0 $X=1444398 $Y=1225650
X1162 14917 15075 15164 15113 25 26 MXI2X1 $T=1450380 1266490 0 180 $X=1447160 $Y=1262550
X1163 14917 15057 15107 15078 25 26 MXI2X1 $T=1450840 1229590 0 180 $X=1447620 $Y=1225650
X1164 14966 14936 15112 15090 25 26 MXI2X1 $T=1448540 1141030 0 0 $X=1448538 $Y=1140778
X1165 12589 475 15153 15226 25 26 MXI2X1 $T=1448540 1185310 1 0 $X=1448538 $Y=1181370
X1166 14867 15247 15200 15115 25 26 MXI2X1 $T=1452680 1118890 0 180 $X=1449460 $Y=1114950
X1167 13390 475 15237 15210 25 26 MXI2X1 $T=1450380 1266490 0 0 $X=1450378 $Y=1266238
X1168 14879 15131 15199 15248 25 26 MXI2X1 $T=1450840 1229590 1 0 $X=1450838 $Y=1225650
X1169 14917 15253 15222 15154 25 26 MXI2X1 $T=1455900 1244350 0 180 $X=1452680 $Y=1240410
X1170 14937 506 15114 15068 25 26 MXI2X1 $T=1456360 1281250 1 180 $X=1453140 $Y=1280998
X1171 14966 14921 15283 15272 25 26 MXI2X1 $T=1454980 1155790 0 0 $X=1454978 $Y=1155538
X1172 14867 15253 15167 15062 25 26 MXI2X1 $T=1458200 1111510 1 180 $X=1454980 $Y=1111258
X1173 14913 15253 15111 15201 25 26 MXI2X1 $T=1458200 1141030 1 180 $X=1454980 $Y=1140778
X1174 497 506 15245 505 25 26 MXI2X1 $T=1458200 1347670 0 180 $X=1454980 $Y=1343730
X1175 14955 15247 15270 15273 25 26 MXI2X1 $T=1455900 1200070 1 0 $X=1455898 $Y=1196130
X1176 13329 475 15257 15314 25 26 MXI2X1 $T=1455900 1266490 0 0 $X=1455898 $Y=1266238
X1177 14879 15296 15263 15262 25 26 MXI2X1 $T=1460040 1207450 0 180 $X=1456820 $Y=1203510
X1178 14913 15131 15343 15260 25 26 MXI2X1 $T=1457280 1126270 0 0 $X=1457278 $Y=1126018
X1179 14926 496 15286 15197 25 26 MXI2X1 $T=1457280 1332910 1 0 $X=1457278 $Y=1328970
X1180 14867 15313 15275 15267 25 26 MXI2X1 $T=1460500 1177930 1 180 $X=1457280 $Y=1177678
X1181 14937 514 15277 15249 25 26 MXI2X1 $T=1460500 1281250 0 180 $X=1457280 $Y=1277310
X1182 15022 496 15212 15118 25 26 MXI2X1 $T=1460500 1296010 1 180 $X=1457280 $Y=1295758
X1183 14913 15313 15294 15244 25 26 MXI2X1 $T=1462340 1155790 1 180 $X=1459120 $Y=1155538
X1184 14966 15253 15323 15291 25 26 MXI2X1 $T=1463720 1118890 0 180 $X=1460500 $Y=1114950
X1185 14913 15352 15337 15274 25 26 MXI2X1 $T=1466020 1148410 0 180 $X=1462800 $Y=1144470
X1186 14955 15313 15338 15373 25 26 MXI2X1 $T=1463260 1192690 1 0 $X=1463258 $Y=1188750
X1187 14926 520 15341 15036 25 26 MXI2X1 $T=1466480 1318150 1 180 $X=1463260 $Y=1317898
X1188 14937 520 15351 15285 25 26 MXI2X1 $T=1468320 1296010 1 180 $X=1465100 $Y=1295758
X1189 14937 517 15332 15369 25 26 MXI2X1 $T=1466020 1281250 1 0 $X=1466018 $Y=1277310
X1190 14867 15131 15346 15214 25 26 MXI2X1 $T=1469240 1126270 1 180 $X=1466020 $Y=1126018
X1191 14867 15296 15359 15316 25 26 MXI2X1 $T=1469240 1177930 1 180 $X=1466020 $Y=1177678
X1192 14929 496 15362 15298 25 26 MXI2X1 $T=1469240 1332910 0 180 $X=1466020 $Y=1328970
X1193 14879 15253 15279 15370 25 26 MXI2X1 $T=1466480 1229590 0 0 $X=1466478 $Y=1229338
X1194 14917 15131 15366 15258 25 26 MXI2X1 $T=1470160 1236970 1 180 $X=1466940 $Y=1236718
X1195 14879 15313 15408 15329 25 26 MXI2X1 $T=1467400 1214830 0 0 $X=1467398 $Y=1214578
X1196 14879 15247 15378 15289 25 26 MXI2X1 $T=1467400 1229590 1 0 $X=1467398 $Y=1225650
X1197 14913 15296 15345 15238 25 26 MXI2X1 $T=1470620 1170550 0 180 $X=1467400 $Y=1166610
X1198 14913 15247 15364 15278 25 26 MXI2X1 $T=1471080 1141030 0 180 $X=1467860 $Y=1137090
X1199 14917 15352 15380 15242 25 26 MXI2X1 $T=1471540 1273870 0 180 $X=1468320 $Y=1269930
X1200 14926 518 15349 15254 25 26 MXI2X1 $T=1471540 1303390 1 180 $X=1468320 $Y=1303138
X1201 497 514 15381 15147 25 26 MXI2X1 $T=1471540 1347670 0 180 $X=1468320 $Y=1343730
X1202 14955 15253 15365 15145 25 26 MXI2X1 $T=1472460 1185310 1 180 $X=1469240 $Y=1185058
X1203 14955 15296 15401 15324 25 26 MXI2X1 $T=1472460 1207450 1 180 $X=1469240 $Y=1207198
X1204 14917 15247 15276 15371 25 26 MXI2X1 $T=1472460 1251730 1 180 $X=1469240 $Y=1251478
X1205 15053 14936 15422 15440 25 26 MXI2X1 $T=1471540 1259110 1 0 $X=1471538 $Y=1255170
X1206 14917 15439 15410 15331 25 26 MXI2X1 $T=1474760 1244350 1 180 $X=1471540 $Y=1244098
X1207 15224 14936 15429 15449 25 26 MXI2X1 $T=1472000 1281250 1 0 $X=1471998 $Y=1277310
X1208 15022 518 15415 15350 25 26 MXI2X1 $T=1475220 1303390 0 180 $X=1472000 $Y=1299450
X1209 14966 15057 15417 15453 25 26 MXI2X1 $T=1472460 1118890 0 0 $X=1472458 $Y=1118638
X1210 15020 14936 15436 15413 25 26 MXI2X1 $T=1472460 1141030 0 0 $X=1472458 $Y=1140778
X1211 14917 15296 15460 15423 25 26 MXI2X1 $T=1472460 1273870 1 0 $X=1472458 $Y=1269930
X1212 497 518 15445 15434 25 26 MXI2X1 $T=1472460 1347670 1 0 $X=1472458 $Y=1343730
X1213 14926 526 15342 15416 25 26 MXI2X1 $T=1475680 1332910 1 180 $X=1472460 $Y=1332658
X1214 15427 14936 15451 15476 25 26 MXI2X1 $T=1472920 1244350 1 0 $X=1472918 $Y=1240410
X1215 14992 15131 15475 15398 25 26 MXI2X1 $T=1473380 1133650 1 0 $X=1473378 $Y=1129710
X1216 14966 15075 15446 15405 25 26 MXI2X1 $T=1473380 1148410 0 0 $X=1473378 $Y=1148158
X1217 14926 517 15461 15477 25 26 MXI2X1 $T=1473380 1332910 1 0 $X=1473378 $Y=1328970
X1218 14913 15439 15430 15424 25 26 MXI2X1 $T=1476600 1155790 1 180 $X=1473380 $Y=1155538
X1219 14993 14921 15431 15420 25 26 MXI2X1 $T=1476600 1185310 0 180 $X=1473380 $Y=1181370
X1220 14917 15313 15414 15335 25 26 MXI2X1 $T=1476600 1266490 0 180 $X=1473380 $Y=1262550
X1221 14992 15057 15403 15399 25 26 MXI2X1 $T=1477060 1141030 0 180 $X=1473840 $Y=1137090
X1222 14926 514 15412 15334 25 26 MXI2X1 $T=1477060 1310770 1 180 $X=1473840 $Y=1310518
X1223 15053 14921 15459 15541 25 26 MXI2X1 $T=1474300 1251730 1 0 $X=1474298 $Y=1247790
X1224 14867 15439 15382 15295 25 26 MXI2X1 $T=1477980 1177930 1 180 $X=1474760 $Y=1177678
X1225 14879 15352 15454 15255 25 26 MXI2X1 $T=1477980 1214830 1 180 $X=1474760 $Y=1214578
X1226 14937 526 15457 15243 25 26 MXI2X1 $T=1478440 1303390 0 180 $X=1475220 $Y=1299450
X1227 14966 15247 15438 15320 25 26 MXI2X1 $T=1475680 1111510 0 0 $X=1475678 $Y=1111258
X1228 13332 475 15426 15455 25 26 MXI2X1 $T=1478900 1222210 1 180 $X=1475680 $Y=1221958
X1229 14929 514 15467 15485 25 26 MXI2X1 $T=1476140 1332910 0 0 $X=1476138 $Y=1332658
X1230 14993 14936 15465 15400 25 26 MXI2X1 $T=1479360 1192690 0 180 $X=1476140 $Y=1188750
X1231 14992 14921 15425 15486 25 26 MXI2X1 $T=1476600 1170550 1 0 $X=1476598 $Y=1166610
X1232 14937 518 15441 15524 25 26 MXI2X1 $T=1479820 1288630 0 0 $X=1479818 $Y=1288378
X1233 14993 15253 15536 15428 25 26 MXI2X1 $T=1480280 1118890 1 0 $X=1480278 $Y=1114950
X1234 14992 14936 15404 15384 25 26 MXI2X1 $T=1486260 1177930 1 180 $X=1483040 $Y=1177678
X1235 14955 15352 15529 15471 25 26 MXI2X1 $T=1486260 1207450 1 180 $X=1483040 $Y=1207198
X1236 15523 14936 15443 15421 25 26 MXI2X1 $T=1486260 1214830 1 180 $X=1483040 $Y=1214578
X1237 14992 15253 15530 15468 25 26 MXI2X1 $T=1486720 1126270 0 180 $X=1483500 $Y=1122330
X1238 14926 506 15507 15406 25 26 MXI2X1 $T=1486720 1303390 1 180 $X=1483500 $Y=1303138
X1239 14879 15439 15540 15458 25 26 MXI2X1 $T=1487640 1200070 1 180 $X=1484420 $Y=1199818
X1240 15022 506 15533 15509 25 26 MXI2X1 $T=1487640 1318150 1 180 $X=1484420 $Y=1317898
X1241 14867 15352 15543 15508 25 26 MXI2X1 $T=1488100 1170550 1 180 $X=1484880 $Y=1170298
X1242 15224 14921 15473 15556 25 26 MXI2X1 $T=1485340 1273870 0 0 $X=1485338 $Y=1273618
X1243 497 520 15546 15472 25 26 MXI2X1 $T=1489020 1347670 1 180 $X=1485800 $Y=1347418
X1244 15022 514 15452 15538 25 26 MXI2X1 $T=1486720 1303390 0 0 $X=1486718 $Y=1303138
X1245 15523 14921 15565 15462 25 26 MXI2X1 $T=1487640 1236970 0 0 $X=1487638 $Y=1236718
X1246 15053 15253 15613 15572 25 26 MXI2X1 $T=1489020 1273870 1 0 $X=1489018 $Y=1269930
X1247 14937 533 15608 15479 25 26 MXI2X1 $T=1489020 1296010 1 0 $X=1489018 $Y=1292070
X1248 15020 15253 15595 15616 25 26 MXI2X1 $T=1489480 1118890 1 0 $X=1489478 $Y=1114950
X1249 15053 15075 15596 15602 25 26 MXI2X1 $T=1489480 1259110 0 0 $X=1489478 $Y=1258858
X1250 14929 506 15621 15525 25 26 MXI2X1 $T=1489480 1340290 0 0 $X=1489478 $Y=1340038
X1251 14993 15075 15567 15549 25 26 MXI2X1 $T=1492700 1200070 1 180 $X=1489480 $Y=1199818
X1252 14926 529 15566 15489 25 26 MXI2X1 $T=1492700 1318150 1 180 $X=1489480 $Y=1317898
X1253 14992 15247 15620 15474 25 26 MXI2X1 $T=1490400 1133650 1 0 $X=1490398 $Y=1129710
X1254 14992 15075 15561 15627 25 26 MXI2X1 $T=1490400 1148410 0 0 $X=1490398 $Y=1148158
X1255 15523 15253 15518 15550 25 26 MXI2X1 $T=1490400 1207450 0 0 $X=1490398 $Y=1207198
X1256 15523 15075 15575 15512 25 26 MXI2X1 $T=1493620 1214830 1 180 $X=1490400 $Y=1214578
X1257 15020 15075 15646 15574 25 26 MXI2X1 $T=1490860 1148410 1 0 $X=1490858 $Y=1144470
X1258 15020 14921 15490 15557 25 26 MXI2X1 $T=1494080 1163170 0 180 $X=1490860 $Y=1159230
X1259 15427 14921 15634 15604 25 26 MXI2X1 $T=1491780 1251730 1 0 $X=1491778 $Y=1247790
X1260 15224 15075 15599 15617 25 26 MXI2X1 $T=1492240 1288630 1 0 $X=1492238 $Y=1284690
X1261 15020 15439 15647 15600 25 26 MXI2X1 $T=1493620 1163170 0 0 $X=1493618 $Y=1162918
X1262 14955 15439 15711 15601 25 26 MXI2X1 $T=1496380 1207450 0 0 $X=1496378 $Y=1207198
X1263 14926 533 15712 15645 25 26 MXI2X1 $T=1503280 1318150 0 180 $X=1500060 $Y=1314210
X1264 15020 15247 15690 15570 25 26 MXI2X1 $T=1503740 1111510 1 180 $X=1500520 $Y=1111258
X1265 15053 15247 15638 15694 25 26 MXI2X1 $T=1503740 1251730 0 180 $X=1500520 $Y=1247790
X1266 15523 15247 15733 15637 25 26 MXI2X1 $T=1505120 1207450 1 180 $X=1501900 $Y=1207198
X1267 15022 520 15554 15662 25 26 MXI2X1 $T=1505580 1296010 1 180 $X=1502360 $Y=1295758
X1268 14929 520 15577 15696 25 26 MXI2X1 $T=1506040 1347670 0 180 $X=1502820 $Y=1343730
X1269 15020 15131 15801 15808 25 26 MXI2X1 $T=1506960 1133650 1 0 $X=1506958 $Y=1129710
X1270 15020 15313 15786 15857 25 26 MXI2X1 $T=1506960 1177930 0 0 $X=1506958 $Y=1177678
X1271 15523 15057 15787 15795 25 26 MXI2X1 $T=1506960 1207450 1 0 $X=1506958 $Y=1203510
X1272 15523 15131 15788 15671 25 26 MXI2X1 $T=1506960 1214830 0 0 $X=1506958 $Y=1214578
X1273 15053 15057 15649 15720 25 26 MXI2X1 $T=1510180 1251730 1 180 $X=1506960 $Y=1251478
X1274 15224 15131 15798 15849 25 26 MXI2X1 $T=1507880 1288630 1 0 $X=1507878 $Y=1284690
X1275 14992 15439 15785 15762 25 26 MXI2X1 $T=1511100 1170550 1 180 $X=1507880 $Y=1170298
X1276 15427 15131 15802 15840 25 26 MXI2X1 $T=1508340 1222210 1 0 $X=1508338 $Y=1218270
X1277 15427 15247 15779 15848 25 26 MXI2X1 $T=1508340 1236970 0 0 $X=1508338 $Y=1236718
X1278 15022 526 15681 15737 25 26 MXI2X1 $T=1511560 1296010 1 180 $X=1508340 $Y=1295758
X1279 15022 533 15794 15746 25 26 MXI2X1 $T=1511560 1318150 1 180 $X=1508340 $Y=1317898
X1280 14993 15247 15846 15745 25 26 MXI2X1 $T=1508800 1118890 1 0 $X=1508798 $Y=1114950
X1281 14993 15131 15832 15777 25 26 MXI2X1 $T=1508800 1141030 1 0 $X=1508798 $Y=1137090
X1282 14992 15352 15797 15853 25 26 MXI2X1 $T=1509260 1148410 1 0 $X=1509258 $Y=1144470
X1283 15053 15131 15812 15639 25 26 MXI2X1 $T=1509260 1251730 1 0 $X=1509258 $Y=1247790
X1284 15020 15296 15659 15767 25 26 MXI2X1 $T=1512480 1163170 1 180 $X=1509260 $Y=1162918
X1285 15224 15247 15650 15607 25 26 MXI2X1 $T=1512480 1273870 1 180 $X=1509260 $Y=1273618
X1286 14929 526 15656 15619 25 26 MXI2X1 $T=1511560 1325530 1 0 $X=1511558 $Y=1321590
X1287 14929 517 15886 15829 25 26 MXI2X1 $T=1513400 1347670 1 0 $X=1513398 $Y=1343730
X1288 15022 517 15878 15796 25 26 MXI2X1 $T=1516620 1310770 0 0 $X=1516618 $Y=1310518
X1289 14966 15313 15844 15896 25 26 MXI2X1 $T=1517540 1163170 0 0 $X=1517538 $Y=1162918
X1290 14993 15296 15929 15856 25 26 MXI2X1 $T=1517540 1192690 0 0 $X=1517538 $Y=1192438
X1291 15020 15352 15876 15793 25 26 MXI2X1 $T=1520760 1148410 0 180 $X=1517540 $Y=1144470
X1292 14993 15439 15877 15834 25 26 MXI2X1 $T=1520760 1200070 1 180 $X=1517540 $Y=1199818
X1293 15427 15313 15783 15774 25 26 MXI2X1 $T=1520760 1251730 0 180 $X=1517540 $Y=1247790
X1294 15224 15057 15854 15749 25 26 MXI2X1 $T=1520760 1273870 1 180 $X=1517540 $Y=1273618
X1295 14929 529 15870 15782 25 26 MXI2X1 $T=1520760 1332910 1 180 $X=1517540 $Y=1332658
X1296 15053 15313 15843 15901 25 26 MXI2X1 $T=1518460 1259110 1 0 $X=1518458 $Y=1255170
X1297 14993 15352 15890 15833 25 26 MXI2X1 $T=1518920 1185310 0 0 $X=1518918 $Y=1185058
X1298 15022 529 15891 15828 25 26 MXI2X1 $T=1518920 1303390 0 0 $X=1518918 $Y=1303138
X1299 14929 533 15902 15841 25 26 MXI2X1 $T=1518920 1325530 0 0 $X=1518918 $Y=1325278
X1300 14992 15296 15961 15956 25 26 MXI2X1 $T=1523520 1185310 0 0 $X=1523518 $Y=1185058
X1301 14993 15057 15920 15847 25 26 MXI2X1 $T=1527200 1141030 0 180 $X=1523980 $Y=1137090
X1302 15523 15439 15900 15719 25 26 MXI2X1 $T=1527200 1214830 0 180 $X=1523980 $Y=1210890
X1303 15523 15352 15979 15987 25 26 MXI2X1 $T=1524900 1229590 1 0 $X=1524898 $Y=1225650
X1304 15523 15313 15999 15976 25 26 MXI2X1 $T=1524900 1251730 1 0 $X=1524898 $Y=1247790
X1305 15224 15313 15970 15874 25 26 MXI2X1 $T=1524900 1288630 0 0 $X=1524898 $Y=1288378
X1306 14926 556 15963 15940 25 26 MXI2X1 $T=1524900 1318150 0 0 $X=1524898 $Y=1317898
X1307 15523 15296 16010 15954 25 26 MXI2X1 $T=1525360 1214830 0 0 $X=1525358 $Y=1214578
X1308 14926 557 15950 15943 25 26 MXI2X1 $T=1525360 1303390 0 0 $X=1525358 $Y=1303138
X1309 14929 557 15958 16012 25 26 MXI2X1 $T=1525360 1325530 1 0 $X=1525358 $Y=1321590
X1310 14966 15352 15951 15931 25 26 MXI2X1 $T=1528580 1148410 0 180 $X=1525360 $Y=1144470
X1311 14966 15439 15930 15855 25 26 MXI2X1 $T=1528580 1155790 1 180 $X=1525360 $Y=1155538
X1312 15053 15439 15892 15827 25 26 MXI2X1 $T=1528580 1259110 0 180 $X=1525360 $Y=1255170
X1313 15224 15296 15957 15813 25 26 MXI2X1 $T=1529040 1273870 1 180 $X=1525820 $Y=1273618
X1314 14966 15296 15948 16049 25 26 MXI2X1 $T=1526740 1163170 0 0 $X=1526738 $Y=1162918
X1315 14955 559 15953 16052 25 26 MXI2X1 $T=1526740 1207450 1 0 $X=1526738 $Y=1203510
X1316 15427 15352 15975 16041 25 26 MXI2X1 $T=1526740 1244350 1 0 $X=1526738 $Y=1240410
X1317 15427 15057 15899 15839 25 26 MXI2X1 $T=1529960 1207450 1 180 $X=1526740 $Y=1207198
X1318 15427 15296 15969 15964 25 26 MXI2X1 $T=1529960 1236970 0 180 $X=1526740 $Y=1233030
X1319 15053 15296 15972 15962 25 26 MXI2X1 $T=1529960 1266490 1 180 $X=1526740 $Y=1266238
X1320 14937 557 15946 15967 25 26 MXI2X1 $T=1529960 1303390 0 180 $X=1526740 $Y=1299450
X1321 14929 556 15988 16005 25 26 MXI2X1 $T=1527200 1340290 1 0 $X=1527198 $Y=1336350
X1322 15224 15439 15966 16054 25 26 MXI2X1 $T=1530880 1288630 0 0 $X=1530878 $Y=1288378
X1323 16008 521 15932 16039 25 26 MXI2X1 $T=1530880 1318150 0 0 $X=1530878 $Y=1317898
X1324 14992 559 16009 15873 25 26 MXI2X1 $T=1534100 1170550 1 180 $X=1530880 $Y=1170298
X1325 15020 15057 15898 15835 25 26 MXI2X1 $T=1531800 1126270 0 0 $X=1531798 $Y=1126018
X1326 15053 15352 16037 15897 25 26 MXI2X1 $T=1531800 1273870 0 0 $X=1531798 $Y=1273618
X1327 14879 559 16031 15916 25 26 MXI2X1 $T=1535020 1214830 1 180 $X=1531800 $Y=1214578
X1328 16027 561 16046 563 25 26 MXI2X1 $T=1532720 1347670 0 0 $X=1532718 $Y=1347418
X1329 15224 15352 16053 15965 25 26 MXI2X1 $T=1534100 1281250 1 0 $X=1534098 $Y=1277310
X1330 14993 559 16058 15982 25 26 MXI2X1 $T=1539160 1200070 0 180 $X=1535940 $Y=1196130
X1331 14937 556 16091 16112 25 26 MXI2X1 $T=1536400 1288630 0 0 $X=1536398 $Y=1288378
X1332 16088 561 16063 16039 25 26 MXI2X1 $T=1539620 1318150 1 180 $X=1536400 $Y=1317898
X1333 14913 559 15936 15872 25 26 MXI2X1 $T=1541000 1141030 1 180 $X=1537780 $Y=1140778
X1334 569 557 16129 16006 25 26 MXI2X1 $T=1540080 1347670 0 0 $X=1540078 $Y=1347418
X1335 14966 559 16097 15994 25 26 MXI2X1 $T=1544220 1148410 0 180 $X=1541000 $Y=1144470
X1336 16172 572 16128 16119 25 26 MXI2X1 $T=1544220 1296010 1 180 $X=1541000 $Y=1295758
X1337 16170 576 15971 16124 25 26 MXI2X1 $T=1544680 1200070 0 180 $X=1541460 $Y=1196130
X1338 15427 559 16007 16103 25 26 MXI2X1 $T=1544680 1222210 1 180 $X=1541460 $Y=1221958
X1339 16178 572 15995 16125 25 26 MXI2X1 $T=1544680 1259110 0 180 $X=1541460 $Y=1255170
X1340 16164 16095 16122 16205 25 26 MXI2X1 $T=1542380 1185310 1 0 $X=1542378 $Y=1181370
X1341 15022 556 16182 15947 25 26 MXI2X1 $T=1542380 1310770 0 0 $X=1542378 $Y=1310518
X1342 16170 572 16149 16231 25 26 MXI2X1 $T=1542840 1185310 0 0 $X=1542838 $Y=1185058
X1343 16171 16095 16150 16202 25 26 MXI2X1 $T=1542840 1207450 0 0 $X=1542838 $Y=1207198
X1344 15053 559 16114 16253 25 26 MXI2X1 $T=1542840 1281250 1 0 $X=1542838 $Y=1277310
X1345 16174 561 16153 16206 25 26 MXI2X1 $T=1542840 1332910 0 0 $X=1542838 $Y=1332658
X1346 16172 576 15804 16221 25 26 MXI2X1 $T=1544220 1296010 0 0 $X=1544218 $Y=1295758
X1347 16211 16095 16084 16183 25 26 MXI2X1 $T=1547440 1177930 0 180 $X=1544220 $Y=1173990
X1348 16183 572 16218 16252 25 26 MXI2X1 $T=1545140 1170550 0 0 $X=1545138 $Y=1170298
X1349 14867 559 16200 16102 25 26 MXI2X1 $T=1548360 1141030 0 180 $X=1545140 $Y=1137090
X1350 16205 572 15960 16228 25 26 MXI2X1 $T=1545600 1177930 0 0 $X=1545598 $Y=1177678
X1351 15523 559 16207 16004 25 26 MXI2X1 $T=1548820 1236970 1 180 $X=1545600 $Y=1236718
X1352 14992 16189 16227 16098 25 26 MXI2X1 $T=1547440 1163170 1 0 $X=1547438 $Y=1159230
X1353 16206 576 16057 16273 25 26 MXI2X1 $T=1547440 1332910 1 0 $X=1547438 $Y=1328970
X1354 15022 557 16173 16283 25 26 MXI2X1 $T=1547900 1310770 0 0 $X=1547898 $Y=1310518
X1355 16249 567 16184 16287 25 26 MXI2X1 $T=1548820 1185310 1 0 $X=1548818 $Y=1181370
X1356 14917 559 16250 16318 25 26 MXI2X1 $T=1550200 1251730 0 0 $X=1550198 $Y=1251478
X1357 14993 16189 16317 16212 25 26 MXI2X1 $T=1552040 1192690 0 0 $X=1552038 $Y=1192438
X1358 14955 16189 16324 16222 25 26 MXI2X1 $T=1552040 1207450 1 0 $X=1552038 $Y=1203510
X1359 14917 16189 16312 16214 25 26 MXI2X1 $T=1552040 1266490 1 0 $X=1552038 $Y=1262550
X1360 16302 564 16194 16280 25 26 MXI2X1 $T=1555260 1244350 1 180 $X=1552040 $Y=1244098
X1361 14879 16189 16220 16325 25 26 MXI2X1 $T=1553420 1214830 0 0 $X=1553418 $Y=1214578
X1362 16298 567 16285 16347 25 26 MXI2X1 $T=1553420 1303390 0 0 $X=1553418 $Y=1303138
X1363 14966 16189 16367 16230 25 26 MXI2X1 $T=1553880 1163170 1 0 $X=1553878 $Y=1159230
X1364 16288 567 16247 16202 25 26 MXI2X1 $T=1553880 1200070 0 0 $X=1553878 $Y=1199818
X1365 16301 567 16248 16345 25 26 MXI2X1 $T=1553880 1214830 1 0 $X=1553878 $Y=1210890
X1366 16299 16095 591 16344 25 26 MXI2X1 $T=1553880 1340290 1 0 $X=1553878 $Y=1336350
X1367 16319 561 16274 16280 25 26 MXI2X1 $T=1557100 1251730 0 180 $X=1553880 $Y=1247790
X1368 16320 572 16160 16297 25 26 MXI2X1 $T=1557100 1273870 0 180 $X=1553880 $Y=1269930
X1369 16304 16095 16294 16333 25 26 MXI2X1 $T=1554340 1236970 1 0 $X=1554338 $Y=1233030
X1370 16307 567 16193 16333 25 26 MXI2X1 $T=1554340 1236970 0 0 $X=1554338 $Y=1236718
X1371 16308 567 592 16344 25 26 MXI2X1 $T=1554340 1347670 0 0 $X=1554338 $Y=1347418
X1372 16326 16095 15998 16287 25 26 MXI2X1 $T=1557560 1177930 1 180 $X=1554340 $Y=1177678
X1373 15427 16189 16303 16203 25 26 MXI2X1 $T=1558020 1229590 0 180 $X=1554800 $Y=1225650
X1374 15020 559 16305 16191 25 26 MXI2X1 $T=1559400 1148410 0 180 $X=1556180 $Y=1144470
X1375 16348 567 16282 16389 25 26 MXI2X1 $T=1558480 1185310 0 0 $X=1558478 $Y=1185058
X1376 14913 16189 16403 16372 25 26 MXI2X1 $T=1559400 1170550 1 0 $X=1559398 $Y=1166610
X1377 16320 576 16295 16407 25 26 MXI2X1 $T=1559400 1273870 1 0 $X=1559398 $Y=1269930
X1378 16347 576 16038 16395 25 26 MXI2X1 $T=1559400 1303390 0 0 $X=1559398 $Y=1303138
X1379 15053 16189 16370 16433 25 26 MXI2X1 $T=1559860 1266490 0 0 $X=1559858 $Y=1266238
X1380 15020 16189 16374 16420 25 26 MXI2X1 $T=1560320 1177930 0 0 $X=1560318 $Y=1177678
X1381 14867 16189 16424 16463 25 26 MXI2X1 $T=1561240 1170550 0 0 $X=1561238 $Y=1170298
X1382 15224 559 16279 16387 25 26 MXI2X1 $T=1564460 1281250 0 180 $X=1561240 $Y=1277310
X1383 16416 16095 16342 16389 25 26 MXI2X1 $T=1564920 1192690 0 180 $X=1561700 $Y=1188750
X1384 16447 16095 16284 16345 25 26 MXI2X1 $T=1568600 1214830 1 180 $X=1565380 $Y=1214578
X1385 15523 16189 16454 16364 25 26 MXI2X1 $T=1565840 1236970 0 0 $X=1565838 $Y=1236718
X1386 16401 561 16357 16455 25 26 MXI2X1 $T=1565840 1288630 1 0 $X=1565838 $Y=1284690
X1387 16467 16095 16437 16429 25 26 MXI2X1 $T=1570440 1170550 0 0 $X=1570438 $Y=1170298
X1388 15224 16189 16481 16441 25 26 MXI2X1 $T=1570440 1281250 1 0 $X=1570438 $Y=1277310
X1389 16487 564 16346 16455 25 26 MXI2X1 $T=1573660 1288630 1 180 $X=1570440 $Y=1288378
X1390 16489 567 16488 16429 25 26 MXI2X1 $T=1572740 1185310 1 0 $X=1572738 $Y=1181370
X1391 9132 26 9049 25 8864 AND2X2 $T=1081000 1185310 0 180 $X=1079160 $Y=1181370
X1392 9151 26 8948 25 9197 AND2X2 $T=1087900 1229590 1 180 $X=1086060 $Y=1229338
X1393 9275 26 9245 25 9255 AND2X2 $T=1089280 1096750 1 180 $X=1087440 $Y=1096498
X1394 9510 26 9438 25 9345 AND2X2 $T=1101240 1236970 1 180 $X=1099400 $Y=1236718
X1395 9438 26 9375 25 9481 AND2X2 $T=1103080 1229590 1 180 $X=1101240 $Y=1229338
X1396 9540 26 9382 25 9636 AND2X2 $T=1103540 1207450 1 0 $X=1103538 $Y=1203510
X1397 9548 26 9379 25 9545 AND2X2 $T=1104920 1163170 0 0 $X=1104918 $Y=1162918
X1398 9344 26 9382 25 9363 AND2X2 $T=1104920 1222210 0 0 $X=1104918 $Y=1221958
X1399 9643 26 9382 25 9392 AND2X2 $T=1106760 1214830 1 180 $X=1104920 $Y=1214578
X1400 9666 26 9382 25 9624 AND2X2 $T=1113200 1214830 1 0 $X=1113198 $Y=1210890
X1401 9800 26 9382 25 9840 AND2X2 $T=1116420 1214830 0 0 $X=1116418 $Y=1214578
X1402 9575 26 9382 25 9920 AND2X2 $T=1121020 1207450 0 0 $X=1121018 $Y=1207198
X1403 10363 26 10428 25 10523 AND2X2 $T=1144940 1347670 1 0 $X=1144938 $Y=1343730
X1404 11074 26 11081 25 11132 AND2X2 $T=1178980 1347670 1 0 $X=1178978 $Y=1343730
X1405 11588 26 11614 25 11538 AND2X2 $T=1207500 1118890 1 0 $X=1207498 $Y=1114950
X1406 15994 26 16121 25 16155 AND2X2 $T=1541000 1148410 0 0 $X=1540998 $Y=1148158
X1407 8917 8822 25 26 8873 AND2XL $T=1062140 1200070 0 180 $X=1060300 $Y=1196130
X1408 8834 8870 25 26 9007 AND2XL $T=1069040 1200070 1 0 $X=1069038 $Y=1196130
X1409 9061 8880 25 26 8982 AND2XL $T=1071340 1207450 0 180 $X=1069500 $Y=1203510
X1410 9199 9116 25 26 9079 AND2XL $T=1081460 1089370 0 180 $X=1079620 $Y=1085430
X1411 9343 8883 25 26 9360 AND2XL $T=1093420 1214830 1 0 $X=1093418 $Y=1210890
X1412 9341 9379 25 26 9492 AND2XL $T=1094800 1155790 0 0 $X=1094798 $Y=1155538
X1413 9238 8980 25 26 9265 AND2XL $T=1096640 1200070 1 180 $X=1094800 $Y=1199818
X1414 9282 9379 25 26 9539 AND2XL $T=1098940 1155790 1 0 $X=1098938 $Y=1151850
X1415 9345 9417 25 26 9575 AND2XL $T=1101240 1236970 1 0 $X=1101238 $Y=1233030
X1416 9417 9436 25 26 9643 AND2XL $T=1105380 1236970 1 0 $X=1105378 $Y=1233030
X1417 9512 9437 25 26 9502 AND2XL $T=1107220 1200070 0 180 $X=1105380 $Y=1196130
X1418 9375 9436 25 26 9666 AND2XL $T=1110440 1236970 1 0 $X=1110438 $Y=1233030
X1419 8948 9151 25 26 9737 AND2XL $T=1110900 1229590 1 0 $X=1110898 $Y=1225650
X1420 10353 10274 25 26 10495 AND2XL $T=1144480 1296010 0 0 $X=1144478 $Y=1295758
X1421 12500 12463 25 26 12630 AND2XL $T=1255340 1185310 1 0 $X=1255338 $Y=1181370
X1422 12685 12889 25 26 13386 AND2XL $T=1297660 1155790 0 180 $X=1295820 $Y=1151850
X1423 8834 25 8814 8862 26 NAND2X1 $T=1058920 1111510 0 0 $X=1058918 $Y=1111258
X1424 8858 25 8863 8904 26 NAND2X1 $T=1059380 1089370 1 0 $X=1059378 $Y=1085430
X1425 8872 25 8884 8911 26 NAND2X1 $T=1060300 1170550 1 0 $X=1060298 $Y=1166610
X1426 8862 25 8882 8962 26 NAND2X1 $T=1060760 1111510 1 0 $X=1060758 $Y=1107570
X1427 8863 25 8923 9014 26 NAND2X1 $T=1065360 1089370 1 0 $X=1065358 $Y=1085430
X1428 8837 25 8919 8974 26 NAND2X1 $T=1065820 1104130 0 0 $X=1065818 $Y=1103878
X1429 8939 25 9002 9084 26 NAND2X1 $T=1069500 1074610 0 0 $X=1069498 $Y=1074358
X1430 8964 25 8816 8837 26 NAND2X1 $T=1069500 1096750 0 0 $X=1069498 $Y=1096498
X1431 9054 25 9043 8946 26 NAND2X1 $T=1072260 1177930 0 180 $X=1070880 $Y=1173990
X1432 9049 25 9043 8932 26 NAND2X1 $T=1072260 1177930 1 180 $X=1070880 $Y=1177678
X1433 9169 25 9049 8943 26 NAND2X1 $T=1076860 1170550 0 180 $X=1075480 $Y=1166610
X1434 9096 25 9080 8916 26 NAND2X1 $T=1076860 1185310 0 180 $X=1075480 $Y=1181370
X1435 9043 25 9090 9096 26 NAND2X1 $T=1075940 1177930 0 0 $X=1075938 $Y=1177678
X1436 9103 25 9091 9082 26 NAND2X1 $T=1077320 1229590 0 180 $X=1075940 $Y=1225650
X1437 9106 25 9073 9154 26 NAND2X1 $T=1077320 1111510 1 0 $X=1077318 $Y=1107570
X1438 9116 25 9048 9231 26 NAND2X1 $T=1077780 1081990 0 0 $X=1077778 $Y=1081738
X1439 9054 25 9132 8872 26 NAND2X1 $T=1079160 1177930 0 180 $X=1077780 $Y=1173990
X1440 9151 25 8883 9103 26 NAND2X1 $T=1079160 1229590 1 180 $X=1077780 $Y=1229338
X1441 9169 25 9090 8677 26 NAND2X1 $T=1080080 1170550 1 0 $X=1080078 $Y=1166610
X1442 9075 25 9194 9224 26 NAND2X1 $T=1081460 1192690 1 0 $X=1081458 $Y=1188750
X1443 9203 25 9127 9219 26 NAND2X1 $T=1082840 1096750 1 0 $X=1082838 $Y=1092810
X1444 9169 25 9054 9141 26 NAND2X1 $T=1084220 1170550 1 0 $X=1084218 $Y=1166610
X1445 9272 25 9132 8920 26 NAND2X1 $T=1087900 1177930 0 180 $X=1086520 $Y=1173990
X1446 9272 25 9043 8859 26 NAND2X1 $T=1088360 1170550 1 180 $X=1086980 $Y=1170298
X1447 9325 25 9277 9266 26 NAND2X1 $T=1089280 1185310 0 180 $X=1087900 $Y=1181370
X1448 9203 25 9281 9275 26 NAND2X1 $T=1089740 1096750 0 180 $X=1088360 $Y=1092810
X1449 9334 25 9049 9177 26 NAND2X1 $T=1090200 1170550 0 180 $X=1088820 $Y=1166610
X1450 9177 25 9271 9415 26 NAND2X1 $T=1092960 1148410 1 0 $X=1092958 $Y=1144470
X1451 9334 25 9090 8741 26 NAND2X1 $T=1092960 1170550 1 0 $X=1092958 $Y=1166610
X1452 9138 25 8961 9210 26 NAND2X1 $T=1094340 1104130 1 180 $X=1092960 $Y=1103878
X1453 9382 25 9343 9128 26 NAND2X1 $T=1094340 1200070 0 180 $X=1092960 $Y=1196130
X1454 9350 25 9345 9335 26 NAND2X1 $T=1094340 1236970 0 180 $X=1092960 $Y=1233030
X1455 9130 25 9324 9327 26 NAND2X1 $T=1093420 1059850 0 0 $X=1093418 $Y=1059598
X1456 8964 25 8931 9357 26 NAND2X1 $T=1093880 1081990 1 0 $X=1093878 $Y=1078050
X1457 9339 25 9389 9397 26 NAND2X1 $T=1095260 1111510 1 0 $X=1095258 $Y=1107570
X1458 9382 25 9360 9358 26 NAND2X1 $T=1095720 1185310 0 0 $X=1095718 $Y=1185058
X1459 9332 25 9403 9469 26 NAND2X1 $T=1096180 1192690 1 0 $X=1096178 $Y=1188750
X1460 9272 25 9334 9359 26 NAND2X1 $T=1096640 1170550 1 0 $X=1096638 $Y=1166610
X1461 9382 25 9354 9487 26 NAND2X1 $T=1096640 1200070 1 0 $X=1096638 $Y=1196130
X1462 9477 25 9427 9232 26 NAND2X1 $T=1098480 1081990 1 180 $X=1097100 $Y=1081738
X1463 9440 25 9439 9517 26 NAND2X1 $T=1098940 1104130 1 0 $X=1098938 $Y=1100190
X1464 9272 25 9169 9353 26 NAND2X1 $T=1098940 1170550 0 0 $X=1098938 $Y=1170298
X1465 9509 25 8732 9325 26 NAND2X1 $T=1100320 1185310 1 180 $X=1098940 $Y=1185058
X1466 9119 25 9432 9548 26 NAND2X1 $T=1099860 1163170 0 0 $X=1099858 $Y=1162918
X1467 9054 25 9334 9119 26 NAND2X1 $T=1100320 1170550 1 0 $X=1100318 $Y=1166610
X1468 9547 25 9535 9417 26 NAND2X1 $T=1104000 1296010 1 180 $X=1102620 $Y=1295758
X1469 9516 25 9563 9657 26 NAND2X1 $T=1104920 1089370 0 0 $X=1104918 $Y=1089118
X1470 9476 25 9597 9661 26 NAND2X1 $T=1105380 1081990 1 0 $X=1105378 $Y=1078050
X1471 9258 25 9101 9440 26 NAND2X1 $T=1106760 1096750 1 180 $X=1105380 $Y=1096498
X1472 9534 25 9102 9516 26 NAND2X1 $T=1111360 1081990 0 180 $X=1109980 $Y=1078050
X1473 9487 25 9690 9555 26 NAND2X1 $T=1111360 1148410 1 180 $X=1109980 $Y=1148158
X1474 9739 25 9691 9559 26 NAND2X1 $T=1111360 1296010 0 180 $X=1109980 $Y=1292070
X1475 8827 25 9708 9689 26 NAND2X1 $T=1112280 1133650 0 180 $X=1110900 $Y=1129710
X1476 9772 25 9726 9715 26 NAND2X1 $T=1113200 1052470 1 180 $X=1111820 $Y=1052218
X1477 9005 25 9708 9797 26 NAND2X1 $T=1112280 1118890 1 0 $X=1112278 $Y=1114950
X1478 8947 25 9624 9813 26 NAND2X1 $T=1113200 1192690 0 0 $X=1113198 $Y=1192438
X1479 8980 25 9708 9875 26 NAND2X1 $T=1115500 1118890 0 0 $X=1115498 $Y=1118638
X1480 9820 25 9824 9894 26 NAND2X1 $T=1116880 1096750 1 0 $X=1116878 $Y=1092810
X1481 9829 25 9520 9932 26 NAND2X1 $T=1117340 1045090 0 0 $X=1117338 $Y=1044838
X1482 9806 25 9270 9820 26 NAND2X1 $T=1118260 1089370 0 0 $X=1118258 $Y=1089118
X1483 9753 25 9755 9901 26 NAND2X1 $T=1118260 1200070 0 0 $X=1118258 $Y=1199818
X1484 51 25 9504 9951 26 NAND2X1 $T=1122860 1133650 1 0 $X=1122858 $Y=1129710
X1485 9382 25 9420 9991 26 NAND2X1 $T=1122860 1185310 0 0 $X=1122858 $Y=1185058
X1486 10106 25 10042 9777 26 NAND2X1 $T=1128380 1096750 0 180 $X=1127000 $Y=1092810
X1487 9996 25 9504 10064 26 NAND2X1 $T=1127460 1207450 0 0 $X=1127458 $Y=1207198
X1488 85 25 9923 9897 26 NAND2X1 $T=1127460 1266490 1 0 $X=1127458 $Y=1262550
X1489 10136 25 9386 9978 26 NAND2X1 $T=1128840 1081990 1 180 $X=1127460 $Y=1081738
X1490 10139 25 10051 10046 26 NAND2X1 $T=1128840 1288630 0 180 $X=1127460 $Y=1284690
X1491 9978 25 9904 9933 26 NAND2X1 $T=1127920 1089370 1 0 $X=1127918 $Y=1085430
X1492 55 25 9504 10066 26 NAND2X1 $T=1127920 1155790 1 0 $X=1127918 $Y=1151850
X1493 87 25 9504 9969 26 NAND2X1 $T=1129300 1111510 1 180 $X=1127920 $Y=1111258
X1494 9243 25 9708 10197 26 NAND2X1 $T=1129300 1133650 1 0 $X=1129298 $Y=1129710
X1495 56 25 9775 10108 26 NAND2X1 $T=1129300 1133650 0 0 $X=1129298 $Y=1133398
X1496 10166 25 9822 10081 26 NAND2X1 $T=1130680 1318150 0 180 $X=1129300 $Y=1314210
X1497 10052 25 10110 10281 26 NAND2X1 $T=1129760 1296010 1 0 $X=1129758 $Y=1292070
X1498 10051 25 10110 10209 26 NAND2X1 $T=1131140 1288630 0 0 $X=1131138 $Y=1288378
X1499 10228 25 10201 9893 26 NAND2X1 $T=1135280 1045090 0 180 $X=1133900 $Y=1041150
X1500 100 25 9504 10078 26 NAND2X1 $T=1136200 1118890 1 180 $X=1134820 $Y=1118638
X1501 10052 25 10139 10291 26 NAND2X1 $T=1135280 1288630 0 0 $X=1135278 $Y=1288378
X1502 70 25 9775 10284 26 NAND2X1 $T=1140800 1185310 1 180 $X=1139420 $Y=1185058
X1503 9437 25 9708 10411 26 NAND2X1 $T=1139880 1141030 0 0 $X=1139878 $Y=1140778
X1504 45 25 9775 9907 26 NAND2X1 $T=1141260 1192690 0 180 $X=1139880 $Y=1188750
X1505 10229 25 9504 10282 26 NAND2X1 $T=1141720 1192690 1 180 $X=1140340 $Y=1192438
X1506 10106 25 10406 10371 26 NAND2X1 $T=1143560 1096750 0 0 $X=1143558 $Y=1096498
X1507 109 25 9775 10325 26 NAND2X1 $T=1145860 1177930 1 180 $X=1144480 $Y=1177678
X1508 9518 25 9708 10520 26 NAND2X1 $T=1144940 1148410 0 0 $X=1144938 $Y=1148158
X1509 9534 25 9518 10392 26 NAND2X1 $T=1146320 1059850 0 180 $X=1144940 $Y=1055910
X1510 10106 25 10438 10400 26 NAND2X1 $T=1145400 1126270 0 0 $X=1145398 $Y=1126018
X1511 10106 25 10466 10181 26 NAND2X1 $T=1146780 1118890 1 0 $X=1146778 $Y=1114950
X1512 10472 25 10492 10462 26 NAND2X1 $T=1149540 1207450 1 180 $X=1148160 $Y=1207198
X1513 111 25 9504 10467 26 NAND2X1 $T=1151840 1133650 1 180 $X=1150460 $Y=1133398
X1514 10435 25 9708 10610 26 NAND2X1 $T=1151380 1155790 0 0 $X=1151378 $Y=1155538
X1515 117 25 9504 10468 26 NAND2X1 $T=1157360 1141030 0 180 $X=1155980 $Y=1137090
X1516 124 25 9504 10638 26 NAND2X1 $T=1158740 1148410 1 180 $X=1157360 $Y=1148158
X1517 10136 25 10435 10583 26 NAND2X1 $T=1157820 1045090 0 0 $X=1157818 $Y=1044838
X1518 10564 25 10744 10798 26 NAND2X1 $T=1162420 1037710 0 0 $X=1162418 $Y=1037458
X1519 10602 25 9708 10746 26 NAND2X1 $T=1163800 1133650 1 180 $X=1162420 $Y=1133398
X1520 139 25 9504 10831 26 NAND2X1 $T=1168860 1133650 1 180 $X=1167480 $Y=1133398
X1521 143 25 9504 10771 26 NAND2X1 $T=1169780 1163170 0 180 $X=1168400 $Y=1159230
X1522 142 25 10880 146 26 NAND2X1 $T=1171160 1340290 0 0 $X=1171158 $Y=1340038
X1523 10934 25 151 11064 26 NAND2X1 $T=1173920 1332910 1 0 $X=1173918 $Y=1328970
X1524 10472 25 11009 10635 26 NAND2X1 $T=1177140 1251730 1 180 $X=1175760 $Y=1251478
X1525 11064 25 11073 11131 26 NAND2X1 $T=1178520 1332910 1 0 $X=1178518 $Y=1328970
X1526 11053 25 11075 156 26 NAND2X1 $T=1179900 1347670 1 180 $X=1178520 $Y=1347418
X1527 161 25 11072 11166 26 NAND2X1 $T=1184040 1325530 1 0 $X=1184038 $Y=1321590
X1528 11081 25 11189 11254 26 NAND2X1 $T=1184040 1347670 1 0 $X=1184038 $Y=1343730
X1529 11189 25 168 11211 26 NAND2X1 $T=1186340 1347670 0 0 $X=1186338 $Y=1347418
X1530 11166 25 11245 11305 26 NAND2X1 $T=1187260 1325530 0 0 $X=1187258 $Y=1325278
X1531 11297 25 11286 170 26 NAND2X1 $T=1190940 1347670 1 180 $X=1189560 $Y=1347418
X1532 11420 25 11343 11286 26 NAND2X1 $T=1193700 1347670 0 180 $X=1192320 $Y=1343730
X1533 182 25 10879 11385 26 NAND2X1 $T=1197380 1318150 1 180 $X=1196000 $Y=1317898
X1534 10972 25 11430 10174 26 NAND2X1 $T=1198760 1229590 0 180 $X=1197380 $Y=1225650
X1535 181 25 11391 11456 26 NAND2X1 $T=1198760 1347670 1 0 $X=1198758 $Y=1343730
X1536 11385 25 11454 11523 26 NAND2X1 $T=1199220 1340290 1 0 $X=1199218 $Y=1336350
X1537 11556 25 11404 11485 26 NAND2X1 $T=1202440 1081990 0 180 $X=1201060 $Y=1078050
X1538 187 25 10906 11433 26 NAND2X1 $T=1203360 1325530 0 180 $X=1201980 $Y=1321590
X1539 11433 25 11605 11595 26 NAND2X1 $T=1207040 1332910 1 0 $X=1207038 $Y=1328970
X1540 11556 25 11596 11587 26 NAND2X1 $T=1210260 1089370 1 180 $X=1208880 $Y=1089118
X1541 11546 25 11052 11614 26 NAND2X1 $T=1209340 1118890 0 0 $X=1209338 $Y=1118638
X1542 11561 25 9624 11621 26 NAND2X1 $T=1213940 1185310 1 180 $X=1212560 $Y=1185058
X1543 11741 25 11564 200 26 NAND2X1 $T=1213480 1340290 0 0 $X=1213478 $Y=1340038
X1544 11425 25 9624 11887 26 NAND2X1 $T=1215780 1170550 0 0 $X=1215778 $Y=1170298
X1545 11799 25 11818 11869 26 NAND2X1 $T=1215780 1185310 1 0 $X=1215778 $Y=1181370
X1546 11556 25 11808 11690 26 NAND2X1 $T=1217160 1052470 1 180 $X=1215780 $Y=1052218
X1547 11601 25 11816 11630 26 NAND2X1 $T=1217160 1104130 0 180 $X=1215780 $Y=1100190
X1548 11926 25 11147 11765 26 NAND2X1 $T=1219000 1111510 1 180 $X=1217620 $Y=1111258
X1549 11721 25 206 11731 26 NAND2X1 $T=1219000 1325530 1 180 $X=1217620 $Y=1325278
X1550 11556 25 11795 11383 26 NAND2X1 $T=1220380 1081990 0 0 $X=1220378 $Y=1081738
X1551 11901 25 11449 11799 26 NAND2X1 $T=1220380 1177930 1 0 $X=1220378 $Y=1173990
X1552 11770 25 11928 209 26 NAND2X1 $T=1222220 1347670 1 180 $X=1220840 $Y=1347418
X1553 11996 25 11721 11626 26 NAND2X1 $T=1223600 1325530 1 180 $X=1222220 $Y=1325278
X1554 11449 25 9708 12007 26 NAND2X1 $T=1223600 1141030 1 0 $X=1223598 $Y=1137090
X1555 11941 25 11437 11601 26 NAND2X1 $T=1225900 1104130 0 180 $X=1224520 $Y=1100190
X1556 211 25 11899 202 26 NAND2X1 $T=1227280 1340290 0 180 $X=1225900 $Y=1336350
X1557 11556 25 12040 11763 26 NAND2X1 $T=1226360 1037710 1 0 $X=1226358 $Y=1033770
X1558 11556 25 11892 12048 26 NAND2X1 $T=1226360 1059850 1 0 $X=1226358 $Y=1055910
X1559 11556 25 11956 12140 26 NAND2X1 $T=1226820 1074610 1 0 $X=1226818 $Y=1070670
X1560 11996 25 192 11992 26 NAND2X1 $T=1226820 1325530 0 0 $X=1226818 $Y=1325278
X1561 220 25 10850 214 26 NAND2X1 $T=1228200 1347670 0 180 $X=1226820 $Y=1343730
X1562 11556 25 12002 11846 26 NAND2X1 $T=1227280 1045090 1 0 $X=1227278 $Y=1041150
X1563 206 25 192 12144 26 NAND2X1 $T=1227740 1332910 1 0 $X=1227738 $Y=1328970
X1564 11314 25 9624 12136 26 NAND2X1 $T=1230960 1163170 1 0 $X=1230958 $Y=1159230
X1565 12141 25 12121 12006 26 NAND2X1 $T=1232340 1104130 0 180 $X=1230960 $Y=1100190
X1566 213 25 9775 11927 26 NAND2X1 $T=1232340 1141030 1 180 $X=1230960 $Y=1140778
X1567 12182 25 12124 12049 26 NAND2X1 $T=1232340 1163170 1 180 $X=1230960 $Y=1162918
X1568 12138 25 10670 12172 26 NAND2X1 $T=1231880 1332910 0 0 $X=1231878 $Y=1332658
X1569 12152 25 12161 12302 26 NAND2X1 $T=1232800 1096750 1 0 $X=1232798 $Y=1092810
X1570 11941 25 11425 12182 26 NAND2X1 $T=1233260 1170550 1 0 $X=1233258 $Y=1166610
X1571 12316 25 12138 12155 26 NAND2X1 $T=1238780 1332910 1 180 $X=1237400 $Y=1332658
X1572 11177 25 9624 12293 26 NAND2X1 $T=1238780 1141030 0 0 $X=1238778 $Y=1140778
X1573 227 25 9775 11751 26 NAND2X1 $T=1241540 1170550 1 180 $X=1240160 $Y=1170298
X1574 10670 25 10729 12358 26 NAND2X1 $T=1242920 1332910 0 0 $X=1242918 $Y=1332658
X1575 12253 25 11322 12141 26 NAND2X1 $T=1243380 1104130 0 0 $X=1243378 $Y=1103878
X1576 11345 25 9624 12304 26 NAND2X1 $T=1244760 1133650 0 180 $X=1243380 $Y=1129710
X1577 12316 25 10729 12352 26 NAND2X1 $T=1243840 1340290 1 0 $X=1243838 $Y=1336350
X1578 231 25 9775 12277 26 NAND2X1 $T=1245220 1155790 1 180 $X=1243840 $Y=1155538
X1579 12391 25 12382 12298 26 NAND2X1 $T=1245220 1163170 0 180 $X=1243840 $Y=1159230
X1580 12463 25 9708 12447 26 NAND2X1 $T=1248900 1148410 1 180 $X=1247520 $Y=1148158
X1581 11220 25 9624 12446 26 NAND2X1 $T=1249820 1155790 0 180 $X=1248440 $Y=1151850
X1582 12545 25 12449 12528 26 NAND2X1 $T=1251660 1052470 1 180 $X=1250280 $Y=1052218
X1583 12594 25 12453 12551 26 NAND2X1 $T=1252580 1067230 1 180 $X=1251200 $Y=1066978
X1584 12604 25 12588 12511 26 NAND2X1 $T=1253500 1074610 0 180 $X=1252120 $Y=1070670
X1585 235 25 9775 12614 26 NAND2X1 $T=1255340 1141030 1 180 $X=1253960 $Y=1140778
X1586 241 25 9775 12495 26 NAND2X1 $T=1255800 1126270 1 180 $X=1254420 $Y=1126018
X1587 242 25 9775 12496 26 NAND2X1 $T=1256260 1141030 0 180 $X=1254880 $Y=1137090
X1588 10972 25 249 12357 26 NAND2X1 $T=1256260 1296010 0 180 $X=1254880 $Y=1292070
X1589 12673 25 12631 12536 26 NAND2X1 $T=1256720 1089370 1 180 $X=1255340 $Y=1089118
X1590 10972 25 254 12587 26 NAND2X1 $T=1260400 1273870 0 180 $X=1259020 $Y=1269930
X1591 10972 25 255 12283 26 NAND2X1 $T=1260400 1281250 0 180 $X=1259020 $Y=1277310
X1592 10972 25 256 12711 26 NAND2X1 $T=1260400 1296010 1 180 $X=1259020 $Y=1295758
X1593 12514 25 9708 12851 26 NAND2X1 $T=1260400 1177930 1 0 $X=1260398 $Y=1173990
X1594 264 25 9504 12764 26 NAND2X1 $T=1266840 1141030 0 180 $X=1265460 $Y=1137090
X1595 12730 25 11225 12604 26 NAND2X1 $T=1267300 1074610 0 180 $X=1265920 $Y=1070670
X1596 12988 25 12829 12539 26 NAND2X1 $T=1267300 1081990 0 180 $X=1265920 $Y=1078050
X1597 12881 25 12849 12756 26 NAND2X1 $T=1267300 1104130 0 180 $X=1265920 $Y=1100190
X1598 12868 25 12916 12910 26 NAND2X1 $T=1266380 1059850 0 0 $X=1266378 $Y=1059598
X1599 12814 25 11344 12673 26 NAND2X1 $T=1267760 1096750 0 0 $X=1267758 $Y=1096498
X1600 10972 25 270 12884 26 NAND2X1 $T=1269140 1251730 1 180 $X=1267760 $Y=1251478
X1601 10972 25 273 12937 26 NAND2X1 $T=1268680 1244350 0 0 $X=1268678 $Y=1244098
X1602 12622 25 9708 13015 26 NAND2X1 $T=1270980 1133650 1 0 $X=1270978 $Y=1129710
X1603 12889 25 9624 13078 26 NAND2X1 $T=1272820 1141030 0 0 $X=1272818 $Y=1140778
X1604 280 25 9504 12890 26 NAND2X1 $T=1274200 1155790 0 180 $X=1272820 $Y=1151850
X1605 12729 25 9624 12931 26 NAND2X1 $T=1274200 1155790 1 180 $X=1272820 $Y=1155538
X1606 279 25 9504 12999 26 NAND2X1 $T=1274200 1177930 0 180 $X=1272820 $Y=1173990
X1607 12927 25 9624 13225 26 NAND2X1 $T=1276960 1133650 0 0 $X=1276958 $Y=1133398
X1608 12874 25 9624 13113 26 NAND2X1 $T=1278340 1170550 0 180 $X=1276960 $Y=1166610
X1609 12582 25 13161 13104 26 NAND2X1 $T=1278340 1059850 1 0 $X=1278338 $Y=1055910
X1610 13232 25 13162 13146 26 NAND2X1 $T=1279720 1067230 1 180 $X=1278340 $Y=1066978
X1611 284 25 9775 13031 26 NAND2X1 $T=1279720 1163170 0 180 $X=1278340 $Y=1159230
X1612 13240 25 13246 13279 26 NAND2X1 $T=1282940 1089370 0 0 $X=1282938 $Y=1089118
X1613 289 25 9775 13117 26 NAND2X1 $T=1284320 1148410 0 180 $X=1282940 $Y=1144470
X1614 12730 25 12926 13261 26 NAND2X1 $T=1283400 1081990 0 0 $X=1283398 $Y=1081738
X1615 300 25 9775 13116 26 NAND2X1 $T=1285240 1133650 0 180 $X=1283860 $Y=1129710
X1616 308 25 9504 13109 26 NAND2X1 $T=1288920 1118890 0 180 $X=1287540 $Y=1114950
X1617 13324 25 13367 13426 26 NAND2X1 $T=1288000 1067230 0 0 $X=1287998 $Y=1066978
X1618 13381 25 13324 13440 26 NAND2X1 $T=1289380 1067230 1 0 $X=1289378 $Y=1063290
X1619 321 25 9504 13127 26 NAND2X1 $T=1290760 1111510 1 180 $X=1289380 $Y=1111258
X1620 12834 25 12729 13418 26 NAND2X1 $T=1289840 1104130 0 0 $X=1289838 $Y=1103878
X1621 309 25 9504 13271 26 NAND2X1 $T=1291680 1133650 1 180 $X=1290300 $Y=1133398
X1622 12253 25 11345 13474 26 NAND2X1 $T=1292140 1118890 1 0 $X=1292138 $Y=1114950
X1623 13361 25 13454 13464 26 NAND2X1 $T=1293520 1089370 0 0 $X=1293518 $Y=1089118
X1624 13459 25 13466 13487 26 NAND2X1 $T=1294440 1104130 1 0 $X=1294438 $Y=1100190
X1625 13499 25 13426 13108 26 NAND2X1 $T=1295820 1052470 1 180 $X=1294440 $Y=1052218
X1626 13240 25 13478 13588 26 NAND2X1 $T=1295820 1096750 1 0 $X=1295818 $Y=1092810
X1627 13427 25 13494 13489 26 NAND2X1 $T=1295820 1133650 0 0 $X=1295818 $Y=1133398
X1628 12154 25 11220 13562 26 NAND2X1 $T=1296740 1148410 1 0 $X=1296738 $Y=1144470
X1629 13488 25 13515 13493 26 NAND2X1 $T=1298120 1118890 0 180 $X=1296740 $Y=1114950
X1630 13651 25 13631 13619 26 NAND2X1 $T=1304100 1118890 1 180 $X=1302720 $Y=1118638
X1631 13418 25 13708 13730 26 NAND2X1 $T=1311920 1104130 1 0 $X=1311918 $Y=1100190
X1632 15804 25 15781 15211 26 NAND2X1 $T=1508800 1296010 0 180 $X=1507420 $Y=1292070
X1633 15932 25 15893 15269 26 NAND2X1 $T=1521680 1318150 1 180 $X=1520300 $Y=1317898
X1634 15971 25 15939 15622 26 NAND2X1 $T=1525820 1192690 1 180 $X=1524440 $Y=1192438
X1635 15960 25 15944 15722 26 NAND2X1 $T=1526280 1177930 1 180 $X=1524900 $Y=1177678
X1636 16038 25 15945 15515 26 NAND2X1 $T=1526280 1310770 0 180 $X=1524900 $Y=1306830
X1637 15998 25 15955 15209 26 NAND2X1 $T=1527200 1155790 0 180 $X=1525820 $Y=1151850
X1638 15995 25 15973 15171 26 NAND2X1 $T=1528580 1251730 1 180 $X=1527200 $Y=1251478
X1639 16057 25 16026 15516 26 NAND2X1 $T=1533180 1332910 0 180 $X=1531800 $Y=1328970
X1640 16075 25 16034 15121 26 NAND2X1 $T=1534100 1259110 0 180 $X=1532720 $Y=1255170
X1641 16046 25 565 15348 26 NAND2X1 $T=1535940 1347670 1 0 $X=1535938 $Y=1343730
X1642 16084 25 16067 15481 26 NAND2X1 $T=1537780 1170550 0 180 $X=1536400 $Y=1166610
X1643 16160 25 16069 15598 26 NAND2X1 $T=1537780 1266490 1 180 $X=1536400 $Y=1266238
X1644 16063 25 16094 15290 26 NAND2X1 $T=1537780 1325530 1 0 $X=1537778 $Y=1321590
X1645 16122 25 16085 15614 26 NAND2X1 $T=1539620 1177930 1 180 $X=1538240 $Y=1177678
X1646 16149 25 16056 15684 26 NAND2X1 $T=1541000 1185310 1 180 $X=1539620 $Y=1185058
X1647 16150 25 16127 15205 26 NAND2X1 $T=1542380 1207450 1 180 $X=1541000 $Y=1207198
X1648 16153 25 16126 15520 26 NAND2X1 $T=1542380 1332910 1 180 $X=1541000 $Y=1332658
X1649 16184 25 16158 15190 26 NAND2X1 $T=1543300 1170550 1 180 $X=1541920 $Y=1170298
X1650 16193 25 16152 15731 26 NAND2X1 $T=1543300 1236970 1 180 $X=1541920 $Y=1236718
X1651 16194 25 16123 15730 26 NAND2X1 $T=1543300 1244350 0 180 $X=1541920 $Y=1240410
X1652 16218 25 16169 15511 26 NAND2X1 $T=1544220 1163170 0 180 $X=1542840 $Y=1159230
X1653 16181 25 16128 15172 26 NAND2X1 $T=1544220 1296010 0 180 $X=1542840 $Y=1292070
X1654 16247 25 16156 15251 26 NAND2X1 $T=1547440 1200070 1 180 $X=1546060 $Y=1199818
X1655 16248 25 16216 15130 26 NAND2X1 $T=1547440 1214830 0 180 $X=1546060 $Y=1210890
X1656 16284 25 16192 15169 26 NAND2X1 $T=1549740 1214830 1 180 $X=1548360 $Y=1214578
X1657 16285 25 16225 15615 26 NAND2X1 $T=1549740 1303390 1 180 $X=1548360 $Y=1303138
X1658 16295 25 16251 15800 26 NAND2X1 $T=1550200 1266490 1 180 $X=1548820 $Y=1266238
X1659 16282 25 16270 15229 26 NAND2X1 $T=1551580 1170550 1 180 $X=1550200 $Y=1170298
X1660 16274 25 16195 15693 26 NAND2X1 $T=1551580 1251730 0 180 $X=1550200 $Y=1247790
X1661 16294 25 16275 15623 26 NAND2X1 $T=1552500 1236970 0 180 $X=1551120 $Y=1233030
X1662 16346 25 16296 15791 26 NAND2X1 $T=1554800 1281250 1 180 $X=1553420 $Y=1280998
X1663 16342 25 16314 15156 26 NAND2X1 $T=1556640 1185310 1 180 $X=1555260 $Y=1185058
X1664 16357 25 16327 15661 26 NAND2X1 $T=1557560 1288630 0 180 $X=1556180 $Y=1284690
X1665 16437 25 16338 15678 26 NAND2X1 $T=1558480 1148410 1 180 $X=1557100 $Y=1148158
X1666 16488 25 16365 15660 26 NAND2X1 $T=1560780 1155790 1 180 $X=1559400 $Y=1155538
X1667 12452 13244 13253 12746 306 13441 13445 25 26 13455 SDFFNSRXL $T=1282480 1281250 1 0 $X=1282478 $Y=1277310
X1668 12313 13280 13299 11826 306 13354 13465 25 26 13557 SDFFNSRXL $T=1284320 1185310 1 0 $X=1284318 $Y=1181370
X1669 12313 13510 13469 11826 306 13354 13280 25 26 13317 SDFFNSRXL $T=1298580 1177930 0 180 $X=1286620 $Y=1173990
X1670 13081 13351 13365 12746 306 13518 13492 25 26 13558 SDFFNSRXL $T=1287080 1303390 0 0 $X=1287078 $Y=1303138
X1671 12452 13314 13375 12746 306 13534 13244 25 26 13561 SDFFNSRXL $T=1287540 1273870 1 0 $X=1287538 $Y=1269930
X1672 13560 13547 13533 11826 320 13374 13363 25 26 13341 SDFFNSRXL $T=1299500 1170550 0 180 $X=1287540 $Y=1166610
X1673 13081 13315 13555 12746 306 13391 13382 25 26 13368 SDFFNSRXL $T=1300420 1332910 1 180 $X=1288460 $Y=1332658
X1674 13560 13363 13347 13599 320 13374 13330 25 26 13460 SDFFNSRXL $T=1306400 1163170 1 180 $X=1294440 $Y=1162918
X1675 13560 13583 13593 11826 336 13690 13547 25 26 13721 SDFFNSRXL $T=1299500 1185310 1 0 $X=1299498 $Y=1181370
X1676 13566 13584 13594 12746 320 13534 13638 25 26 13785 SDFFNSRXL $T=1299500 1273870 1 0 $X=1299498 $Y=1269930
X1677 13560 13589 13598 13599 337 13694 13642 25 26 13720 SDFFNSRXL $T=1299960 1148410 0 0 $X=1299958 $Y=1148158
X1678 13566 13600 13610 12746 338 13707 13388 25 26 13793 SDFFNSRXL $T=1300420 1259110 0 0 $X=1300418 $Y=1258858
X1679 13081 13492 13611 12746 338 13518 13618 25 26 13804 SDFFNSRXL $T=1300420 1303390 0 0 $X=1300418 $Y=1303138
X1680 13560 341 13692 11826 306 13354 13510 25 26 13580 SDFFNSRXL $T=1312380 1177930 1 180 $X=1300420 $Y=1177678
X1681 13560 13607 13614 11826 306 13712 13502 25 26 13723 SDFFNSRXL $T=1300880 1192690 0 0 $X=1300878 $Y=1192438
X1682 13560 13634 13683 13599 320 13374 13606 25 26 13592 SDFFNSRXL $T=1312840 1170550 0 180 $X=1300880 $Y=1166610
X1683 13560 13606 13657 11826 320 13354 13583 25 26 13877 SDFFNSRXL $T=1303180 1177930 1 0 $X=1303178 $Y=1173990
X1684 13081 13601 13648 12746 338 13391 13636 25 26 13749 SDFFNSRXL $T=1303180 1332910 0 0 $X=1303178 $Y=1332658
X1685 13349 13685 13713 13687 320 13660 13650 25 26 13637 SDFFNSRXL $T=1315140 1251730 0 180 $X=1303180 $Y=1247790
X1686 13566 13733 13682 12746 320 13441 13584 25 26 13630 SDFFNSRXL $T=1315140 1281250 1 180 $X=1303180 $Y=1280998
X1687 13640 13656 13666 13599 339 13734 13716 25 26 13753 SDFFNSRXL $T=1303640 1126270 1 0 $X=1303638 $Y=1122330
X1688 13560 13632 13604 13599 320 13694 13589 25 26 13754 SDFFNSRXL $T=1303640 1148410 1 0 $X=1303638 $Y=1144470
X1689 13560 13633 13605 13599 338 13735 13634 25 26 13755 SDFFNSRXL $T=1303640 1163170 1 0 $X=1303638 $Y=1159230
X1690 13081 13658 13664 12746 340 13736 13747 25 26 13761 SDFFNSRXL $T=1303640 1296010 0 0 $X=1303638 $Y=1295758
X1691 13560 13661 13641 13599 320 13671 13632 25 26 13767 SDFFNSRXL $T=1304100 1141030 0 0 $X=1304098 $Y=1140778
X1692 13560 13642 13668 13599 337 13694 13662 25 26 13790 SDFFNSRXL $T=1304100 1155790 1 0 $X=1304098 $Y=1151850
X1693 13560 13662 13643 13599 338 13694 13633 25 26 13780 SDFFNSRXL $T=1304100 1155790 0 0 $X=1304098 $Y=1155538
X1694 13560 13465 13672 11826 306 13712 13607 25 26 13769 SDFFNSRXL $T=1304100 1192690 1 0 $X=1304098 $Y=1188750
X1695 13609 13256 13673 11826 306 13738 13663 25 26 13791 SDFFNSRXL $T=1304100 1207450 1 0 $X=1304098 $Y=1203510
X1696 13081 13638 13674 12746 340 13736 13658 25 26 13807 SDFFNSRXL $T=1304100 1296010 1 0 $X=1304098 $Y=1292070
X1697 13081 13591 13670 12746 338 13518 13693 25 26 13824 SDFFNSRXL $T=1304100 1310770 0 0 $X=1304098 $Y=1310518
X1698 13081 13665 13647 12746 306 13741 13601 25 26 13765 SDFFNSRXL $T=1304100 1332910 1 0 $X=1304098 $Y=1328970
X1699 13640 13716 13719 13599 339 13671 13661 25 26 13654 SDFFNSRXL $T=1316060 1133650 0 180 $X=1304100 $Y=1129710
X1700 348 13743 13724 12746 306 13391 310 25 26 13655 SDFFNSRXL $T=1316060 1340290 0 180 $X=1304100 $Y=1336350
X1701 13349 13608 13645 11826 306 13744 13491 25 26 13783 SDFFNSRXL $T=1304560 1222210 0 0 $X=1304558 $Y=1221958
X1702 13349 13669 13678 11826 338 13745 13685 25 26 13775 SDFFNSRXL $T=1304560 1229590 0 0 $X=1304558 $Y=1229338
X1703 13349 13623 13564 13687 306 13746 13458 25 26 13784 SDFFNSRXL $T=1304560 1244350 1 0 $X=1304558 $Y=1240410
X1704 13081 13603 13680 12746 338 13741 13665 25 26 13788 SDFFNSRXL $T=1304560 1325530 1 0 $X=1304558 $Y=1321590
X1705 13640 13751 13710 13599 342 13677 13656 25 26 13659 SDFFNSRXL $T=1316520 1118890 0 180 $X=1304560 $Y=1114950
X1706 13646 13505 13627 13687 306 13660 13600 25 26 13792 SDFFNSRXL $T=1305020 1251730 0 0 $X=1305018 $Y=1251478
X1707 13349 13686 13688 13687 336 13745 13669 25 26 13819 SDFFNSRXL $T=1307780 1236970 1 0 $X=1307778 $Y=1233030
X1708 13566 13650 13706 13687 340 13660 13826 25 26 13886 SDFFNSRXL $T=1309160 1259110 1 0 $X=1309158 $Y=1255170
X1709 13566 13742 13756 13687 338 13707 13760 25 26 13882 SDFFNSRXL $T=1313760 1266490 1 0 $X=1313758 $Y=1262550
X1710 13609 13752 13759 11826 340 13875 13872 25 26 13887 SDFFNSRXL $T=1314220 1214830 0 0 $X=1314218 $Y=1214578
X1711 13566 13760 13772 12746 336 13441 13771 25 26 13869 SDFFNSRXL $T=1314680 1273870 0 0 $X=1314678 $Y=1273618
X1712 348 13878 13827 12746 337 13518 13762 25 26 13748 SDFFNSRXL $T=1326640 1310770 0 180 $X=1314680 $Y=1306830
X1713 13640 13858 13809 13599 338 13694 13774 25 26 13763 SDFFNSRXL $T=1327560 1148410 0 180 $X=1315600 $Y=1144470
X1714 13560 13774 13802 13599 339 13671 13855 25 26 13944 SDFFNSRXL $T=1316520 1141030 0 0 $X=1316518 $Y=1140778
X1715 13081 13794 13798 12746 337 13741 13850 25 26 13870 SDFFNSRXL $T=1316520 1325530 0 0 $X=1316518 $Y=1325278
X1716 13640 13805 13812 13599 13851 13901 13840 25 26 13907 SDFFNSRXL $T=1317440 1111510 1 0 $X=1317438 $Y=1107570
X1717 13609 13806 13810 11826 320 13744 13742 25 26 13904 SDFFNSRXL $T=1317440 1222210 0 0 $X=1317438 $Y=1221958
X1718 13640 13813 13820 13599 13851 13901 13805 25 26 13914 SDFFNSRXL $T=1318360 1104130 1 0 $X=1318358 $Y=1100190
X1719 13609 13814 13818 11826 340 13738 13752 25 26 13916 SDFFNSRXL $T=1318360 1207450 0 0 $X=1318358 $Y=1207198
X1720 348 13636 13799 12746 338 13890 13743 25 26 383 SDFFNSRXL $T=1318360 1340290 0 0 $X=1318358 $Y=1340038
X1721 13560 13815 13825 11826 336 13690 13908 25 26 13860 SDFFNSRXL $T=1318820 1185310 1 0 $X=1318818 $Y=1181370
X1722 13609 13822 13830 11826 337 13892 13814 25 26 13997 SDFFNSRXL $T=1319280 1207450 1 0 $X=1319278 $Y=1203510
X1723 13349 13821 13829 13687 13851 13745 13686 25 26 13945 SDFFNSRXL $T=1319280 1236970 0 0 $X=1319278 $Y=1236718
X1724 13560 13841 13845 13599 337 13694 13858 25 26 13859 SDFFNSRXL $T=1320200 1155790 0 0 $X=1320198 $Y=1155538
X1725 13566 13930 13848 12746 336 13736 356 25 26 13844 SDFFNSRXL $T=1333080 1288630 0 180 $X=1321120 $Y=1284690
X1726 13640 13840 13854 13599 362 13677 13751 25 26 13995 SDFFNSRXL $T=1321580 1118890 1 0 $X=1321578 $Y=1114950
X1727 348 13850 13862 12746 337 13391 13922 25 26 13871 SDFFNSRXL $T=1321580 1340290 1 0 $X=1321578 $Y=1336350
X1728 13566 13946 13909 12746 337 13518 13849 25 26 13779 SDFFNSRXL $T=1333540 1303390 0 180 $X=1321580 $Y=1299450
X1729 13349 13856 13846 13687 338 13746 13842 25 26 13963 SDFFNSRXL $T=1322040 1244350 1 0 $X=1322038 $Y=1240410
X1730 13349 13842 13864 13687 337 13948 13847 25 26 13905 SDFFNSRXL $T=1322040 1251730 1 0 $X=1322038 $Y=1247790
X1731 13640 13808 13950 13599 362 13677 13857 25 26 13852 SDFFNSRXL $T=1334460 1118890 1 180 $X=1322500 $Y=1118638
X1732 13566 13826 13898 13687 342 13707 13910 25 26 14058 SDFFNSRXL $T=1325720 1266490 1 0 $X=1325718 $Y=1262550
X1733 13609 13872 13899 13687 342 13875 13959 25 26 14009 SDFFNSRXL $T=1326180 1214830 0 0 $X=1326178 $Y=1214578
X1734 348 13900 13861 12746 13851 13518 13878 25 26 14060 SDFFNSRXL $T=1326640 1310770 0 0 $X=1326638 $Y=1310518
X1735 348 14053 14050 12746 390 13924 13900 25 26 13911 SDFFNSRXL $T=1341360 1318150 0 180 $X=1329400 $Y=1314210
X1736 13640 13857 13941 13599 13851 13901 14062 25 26 14087 SDFFNSRXL $T=1330320 1104130 1 0 $X=1330318 $Y=1100190
X1737 13566 14068 13978 13687 13851 13441 13930 25 26 13923 SDFFNSRXL $T=1342740 1273870 1 180 $X=1330780 $Y=1273618
X1738 13942 14094 13996 13599 339 13374 13758 25 26 13947 SDFFNSRXL $T=1344120 1170550 0 180 $X=1332160 $Y=1166610
X1739 13942 13967 13982 13599 13851 13694 13951 25 26 14296 SDFFNSRXL $T=1334000 1155790 0 0 $X=1333998 $Y=1155538
X1740 13349 13970 13917 13687 339 13948 13921 25 26 14035 SDFFNSRXL $T=1334000 1251730 1 0 $X=1333998 $Y=1247790
X1741 348 13874 13990 12746 362 13391 14006 25 26 14120 SDFFNSRXL $T=1334460 1340290 1 0 $X=1334458 $Y=1336350
X1742 13349 14088 14112 13687 342 13746 13970 25 26 13976 SDFFNSRXL $T=1346880 1244350 0 180 $X=1334920 $Y=1240410
X1743 13609 13908 13969 13998 342 13712 13770 25 26 14184 SDFFNSRXL $T=1335380 1192690 1 0 $X=1335378 $Y=1188750
X1744 13609 14092 14113 13687 339 13744 13867 25 26 13983 SDFFNSRXL $T=1347340 1229590 0 180 $X=1335380 $Y=1225650
X1745 13566 14004 14014 12746 339 13441 14005 25 26 14169 SDFFNSRXL $T=1335840 1281250 0 0 $X=1335838 $Y=1280998
X1746 348 14006 14013 12746 362 13391 14020 25 26 14153 SDFFNSRXL $T=1335840 1332910 1 0 $X=1335838 $Y=1328970
X1747 13942 14003 14010 13599 13851 14022 13967 25 26 14001 SDFFNSRXL $T=1348260 1148410 0 180 $X=1336300 $Y=1144470
X1748 13942 14016 14030 13998 362 13712 14029 25 26 14219 SDFFNSRXL $T=1336760 1192690 0 0 $X=1336758 $Y=1192438
X1749 13942 14028 13987 13998 338 13354 14003 25 26 14137 SDFFNSRXL $T=1337220 1177930 1 0 $X=1337218 $Y=1173990
X1750 348 14002 14036 12746 13851 13518 14129 25 26 14142 SDFFNSRXL $T=1337220 1303390 1 0 $X=1337218 $Y=1299450
X1751 392 14032 394 243 390 13890 400 25 26 402 SDFFNSRXL $T=1337220 1347670 0 0 $X=1337218 $Y=1347418
X1752 13609 14041 14043 13998 13851 13892 14016 25 26 14220 SDFFNSRXL $T=1338140 1200070 1 0 $X=1338138 $Y=1196130
X1753 13609 14042 14044 13998 390 13875 14064 25 26 14168 SDFFNSRXL $T=1338140 1214830 0 0 $X=1338138 $Y=1214578
X1754 13566 13910 14049 13687 342 13660 14052 25 26 14093 SDFFNSRXL $T=1338140 1259110 1 0 $X=1338138 $Y=1255170
X1755 13640 14027 14054 13599 342 14136 14148 25 26 14101 SDFFNSRXL $T=1338600 1133650 1 0 $X=1338598 $Y=1129710
X1756 13609 14029 14051 13998 390 13690 14028 25 26 14178 SDFFNSRXL $T=1338600 1185310 0 0 $X=1338598 $Y=1185058
X1757 13609 13959 13999 13687 342 13875 13806 25 26 14210 SDFFNSRXL $T=1338600 1222210 1 0 $X=1338598 $Y=1218270
X1758 348 14045 13980 12746 390 13518 13946 25 26 14061 SDFFNSRXL $T=1338600 1303390 0 0 $X=1338598 $Y=1303138
X1759 348 14046 14056 396 13851 13924 14045 25 26 14154 SDFFNSRXL $T=1338600 1318150 0 0 $X=1338598 $Y=1317898
X1760 13640 14062 13994 13599 362 13901 14024 25 26 14008 SDFFNSRXL $T=1350560 1111510 0 180 $X=1338600 $Y=1107570
X1761 14150 14020 14118 396 13851 13741 14046 25 26 14037 SDFFNSRXL $T=1350560 1325530 1 180 $X=1338600 $Y=1325278
X1762 13566 14052 14012 13687 342 13534 14034 25 26 14172 SDFFNSRXL $T=1339060 1273870 1 0 $X=1339058 $Y=1269930
X1763 13640 14095 14115 13599 362 13901 13813 25 26 14039 SDFFNSRXL $T=1351020 1096750 1 180 $X=1339060 $Y=1096498
X1764 13566 13849 14066 12746 390 14149 14100 25 26 14173 SDFFNSRXL $T=1339520 1288630 1 0 $X=1339518 $Y=1284690
X1765 13609 14064 14084 13998 342 13892 13952 25 26 14190 SDFFNSRXL $T=1340440 1200070 0 0 $X=1340438 $Y=1199818
X1766 13349 14122 14134 13687 362 13746 14092 25 26 14070 SDFFNSRXL $T=1353320 1244350 1 180 $X=1341360 $Y=1244098
X1767 13640 14188 14185 13599 362 13901 14095 25 26 14091 SDFFNSRXL $T=1354240 1104130 0 180 $X=1342280 $Y=1100190
X1768 13566 14034 14105 13687 342 13441 14004 25 26 14206 SDFFNSRXL $T=1342740 1273870 0 0 $X=1342738 $Y=1273618
X1769 13566 14100 14059 396 13851 14195 14090 25 26 14212 SDFFNSRXL $T=1342740 1296010 0 0 $X=1342738 $Y=1295758
X1770 13566 13921 14089 13687 13851 13534 14068 25 26 14103 SDFFNSRXL $T=1343660 1266490 0 0 $X=1343658 $Y=1266238
X1771 348 14129 14133 396 390 14233 14053 25 26 14126 SDFFNSRXL $T=1346420 1318150 1 0 $X=1346418 $Y=1314210
X1772 13349 14130 14117 13687 342 13660 14122 25 26 14250 SDFFNSRXL $T=1346880 1251730 0 0 $X=1346878 $Y=1251478
X1773 13942 14155 14167 13998 362 13374 14234 25 26 14285 SDFFNSRXL $T=1349640 1170550 0 0 $X=1349638 $Y=1170298
X1774 14150 14090 14170 396 13851 14195 14213 25 26 14114 SDFFNSRXL $T=1349640 1303390 1 0 $X=1349638 $Y=1299450
X1775 13609 14267 14263 13998 362 13738 14041 25 26 14145 SDFFNSRXL $T=1361600 1207450 0 180 $X=1349640 $Y=1203510
X1776 13640 14183 14189 13599 406 13677 14269 25 26 14253 SDFFNSRXL $T=1351480 1118890 1 0 $X=1351478 $Y=1114950
X1777 13942 14303 14209 13998 417 13735 14155 25 26 14186 SDFFNSRXL $T=1364360 1163170 1 180 $X=1352400 $Y=1162918
X1778 13349 14249 14193 13687 342 13745 14085 25 26 14176 SDFFNSRXL $T=1364820 1229590 1 180 $X=1352860 $Y=1229338
X1779 13349 14314 14311 13687 390 13707 14204 25 26 14198 SDFFNSRXL $T=1365280 1259110 0 180 $X=1353320 $Y=1255170
X1780 13942 14148 14223 13599 406 14136 14336 25 26 14255 SDFFNSRXL $T=1354240 1133650 1 0 $X=1354238 $Y=1129710
X1781 14284 14323 14304 13599 420 13901 14188 25 26 14201 SDFFNSRXL $T=1366200 1104130 0 180 $X=1354240 $Y=1100190
X1782 13349 14344 14334 13687 13851 13746 14130 25 26 14216 SDFFNSRXL $T=1367120 1244350 0 180 $X=1355160 $Y=1240410
X1783 14150 14349 14106 396 13851 13391 14104 25 26 14182 SDFFNSRXL $T=1367580 1340290 0 180 $X=1355620 $Y=1336350
X1784 13942 14234 14238 13998 13851 13690 14297 25 26 14298 SDFFNSRXL $T=1356080 1185310 1 0 $X=1356078 $Y=1181370
X1785 14465 14364 14362 13687 417 13745 14249 25 26 14239 SDFFNSRXL $T=1369420 1236970 1 180 $X=1357460 $Y=1236718
X1786 14284 14374 14368 13599 406 13677 14183 25 26 14247 SDFFNSRXL $T=1370340 1118890 1 180 $X=1358380 $Y=1118638
X1787 14284 14269 14300 13599 13851 14403 14323 25 26 14208 SDFFNSRXL $T=1361140 1111510 0 0 $X=1361138 $Y=1111258
X1788 14465 14477 14473 13687 417 13534 14345 25 26 14312 SDFFNSRXL $T=1377240 1273870 0 180 $X=1365280 $Y=1269930
X1789 428 14104 14363 396 418 13890 14461 25 26 14446 SDFFNSRXL $T=1366200 1347670 1 0 $X=1366198 $Y=1343730
X1790 13942 14327 14370 13998 406 13738 14267 25 26 14499 SDFFNSRXL $T=1367120 1207450 0 0 $X=1367118 $Y=1207198
X1791 14150 14378 14389 396 438 14502 14455 25 26 14483 SDFFNSRXL $T=1368500 1296010 0 0 $X=1368498 $Y=1295758
X1792 14284 14399 14421 13998 420 13734 14374 25 26 14315 SDFFNSRXL $T=1380460 1126270 1 180 $X=1368500 $Y=1126018
X1793 14150 14442 14504 396 438 14391 14349 25 26 14372 SDFFNSRXL $T=1380460 1332910 0 180 $X=1368500 $Y=1328970
X1794 14400 14508 14506 13998 417 13694 14303 25 26 14301 SDFFNSRXL $T=1380920 1155790 1 180 $X=1368960 $Y=1155538
X1795 14518 14297 14443 13998 438 13354 14381 25 26 14376 SDFFNSRXL $T=1380920 1177930 1 180 $X=1368960 $Y=1177678
X1796 14465 14486 14459 13687 406 13707 14364 25 26 14360 SDFFNSRXL $T=1380920 1259110 0 180 $X=1368960 $Y=1255170
X1797 13942 14397 14396 13998 418 13690 14428 25 26 14453 SDFFNSRXL $T=1369880 1185310 0 0 $X=1369878 $Y=1185058
X1798 14465 14454 14384 13687 420 14405 14344 25 26 14387 SDFFNSRXL $T=1381840 1244350 0 180 $X=1369880 $Y=1240410
X1799 14400 14456 14511 13599 438 13677 14398 25 26 14271 SDFFNSRXL $T=1382300 1118890 1 180 $X=1370340 $Y=1118638
X1800 14150 14338 14423 396 438 14233 14451 25 26 14525 SDFFNSRXL $T=1370800 1318150 1 0 $X=1370798 $Y=1314210
X1801 13942 14422 14343 13998 438 13892 14327 25 26 14556 SDFFNSRXL $T=1371260 1200070 0 0 $X=1371258 $Y=1199818
X1802 14400 14457 14395 13998 438 14136 14399 25 26 14235 SDFFNSRXL $T=1383220 1133650 1 180 $X=1371260 $Y=1133398
X1803 14400 14537 14426 13599 420 13901 14420 25 26 14225 SDFFNSRXL $T=1383680 1096750 1 180 $X=1371720 $Y=1096498
X1804 14400 14425 14462 13599 406 14403 14514 25 26 14540 SDFFNSRXL $T=1373100 1111510 1 0 $X=1373098 $Y=1107570
X1805 13942 14448 14429 13998 418 14544 14422 25 26 14552 SDFFNSRXL $T=1373100 1200070 1 0 $X=1373098 $Y=1196130
X1806 14150 14451 14460 396 418 14546 14442 25 26 14513 SDFFNSRXL $T=1373100 1325530 0 0 $X=1373098 $Y=1325278
X1807 14400 14420 14419 13599 420 13901 14425 25 26 14433 SDFFNSRXL $T=1385060 1104130 1 180 $X=1373100 $Y=1103878
X1808 13942 14548 14545 13998 406 13875 14444 25 26 14436 SDFFNSRXL $T=1385060 1222210 0 180 $X=1373100 $Y=1218270
X1809 14150 14549 14469 13687 418 14466 14314 25 26 14438 SDFFNSRXL $T=1385060 1273870 1 180 $X=1373100 $Y=1273618
X1810 428 14461 439 396 418 444 446 25 26 443 SDFFNSRXL $T=1373560 1347670 0 0 $X=1373558 $Y=1347418
X1811 14400 14514 14522 13599 438 13677 14456 25 26 14440 SDFFNSRXL $T=1385520 1118890 0 180 $X=1373560 $Y=1114950
X1812 14400 14398 14551 13998 438 14136 14457 25 26 14256 SDFFNSRXL $T=1385520 1133650 0 180 $X=1373560 $Y=1129710
X1813 14400 14266 14447 13998 418 13671 14452 25 26 14463 SDFFNSRXL $T=1386440 1141030 0 180 $X=1374480 $Y=1137090
X1814 14400 14487 14492 13998 418 14022 14508 25 26 14595 SDFFNSRXL $T=1376320 1148410 0 0 $X=1376318 $Y=1148158
X1815 14465 14345 14541 13687 438 13707 14486 25 26 14299 SDFFNSRXL $T=1388280 1266490 0 180 $X=1376320 $Y=1262550
X1816 14150 14572 14512 13687 417 13534 14477 25 26 14489 SDFFNSRXL $T=1389200 1273870 0 180 $X=1377240 $Y=1269930
X1817 14465 14204 14509 13687 420 13948 14610 25 26 14632 SDFFNSRXL $T=1378160 1251730 1 0 $X=1378158 $Y=1247790
X1818 14518 14381 14538 13998 420 13690 14448 25 26 14432 SDFFNSRXL $T=1391500 1185310 0 180 $X=1379540 $Y=1181370
X1819 14150 14620 14470 396 438 14195 14378 25 26 14510 SDFFNSRXL $T=1391500 1303390 1 180 $X=1379540 $Y=1303138
X1820 14150 14562 14625 396 420 14149 14519 25 26 14439 SDFFNSRXL $T=1391960 1288630 0 180 $X=1380000 $Y=1284690
X1821 14400 14452 14557 13998 14596 14022 14487 25 26 14638 SDFFNSRXL $T=1383220 1148410 1 0 $X=1383218 $Y=1144470
X1822 14465 14617 14630 13687 438 14580 14569 25 26 14337 SDFFNSRXL $T=1397480 1259110 1 180 $X=1385520 $Y=1258858
X1823 14465 14624 14588 13687 406 14466 14572 25 26 14561 SDFFNSRXL $T=1397480 1273870 1 180 $X=1385520 $Y=1273618
X1824 14400 14573 14583 13599 420 14403 14685 25 26 14700 SDFFNSRXL $T=1385980 1111510 1 0 $X=1385978 $Y=1107570
X1825 13942 14575 14584 13998 406 13712 14615 25 26 14494 SDFFNSRXL $T=1385980 1192690 0 0 $X=1385978 $Y=1192438
X1826 14465 14488 14585 13687 418 13745 14472 25 26 14677 SDFFNSRXL $T=1385980 1236970 0 0 $X=1385978 $Y=1236718
X1827 14518 14682 14609 13998 455 14586 14574 25 26 14567 SDFFNSRXL $T=1397940 1177930 0 180 $X=1385980 $Y=1173990
X1828 14150 14591 14679 396 420 14546 14582 25 26 14503 SDFFNSRXL $T=1397940 1325530 1 180 $X=1385980 $Y=1325278
X1829 14599 14683 14680 396 420 14391 14578 25 26 14491 SDFFNSRXL $T=1397940 1332910 0 180 $X=1385980 $Y=1328970
X1830 14518 14574 14587 13998 455 14586 14397 25 26 14669 SDFFNSRXL $T=1386440 1177930 0 0 $X=1386438 $Y=1177678
X1831 14400 14600 14603 13599 438 14403 14573 25 26 14571 SDFFNSRXL $T=1398400 1111510 1 180 $X=1386440 $Y=1111258
X1832 13942 14592 14605 13998 14596 14691 14696 25 26 14710 SDFFNSRXL $T=1387360 1207450 1 0 $X=1387358 $Y=1203510
X1833 14465 14593 14606 13687 420 14580 14617 25 26 14707 SDFFNSRXL $T=1387360 1259110 1 0 $X=1387358 $Y=1255170
X1834 14400 14685 14694 13599 420 13901 14537 25 26 14579 SDFFNSRXL $T=1399780 1104130 0 180 $X=1387820 $Y=1100190
X1835 14400 14662 14695 13599 438 13906 14600 25 26 14590 SDFFNSRXL $T=1399780 1118890 1 180 $X=1387820 $Y=1118638
X1836 14607 14519 14618 396 455 14149 14676 25 26 14740 SDFFNSRXL $T=1388740 1288630 0 0 $X=1388738 $Y=1288378
X1837 14518 14612 14701 13998 420 14623 14575 25 26 14539 SDFFNSRXL $T=1400700 1192690 0 180 $X=1388740 $Y=1188750
X1838 14599 14621 14631 396 455 14233 14646 25 26 14736 SDFFNSRXL $T=1389200 1318150 1 0 $X=1389198 $Y=1314210
X1839 14732 14706 14670 13998 420 13875 14548 25 26 14394 SDFFNSRXL $T=1401160 1222210 0 180 $X=1389200 $Y=1218270
X1840 14599 462 14602 396 460 444 14613 25 26 449 SDFFNSRXL $T=1401160 1347670 1 180 $X=1389200 $Y=1347418
X1841 14465 14635 14703 13687 438 13744 14593 25 26 14445 SDFFNSRXL $T=1401620 1229590 0 180 $X=1389660 $Y=1225650
X1842 14465 14569 14667 13687 438 13534 14624 25 26 14524 SDFFNSRXL $T=1401620 1273870 0 180 $X=1389660 $Y=1269930
X1843 14150 14626 14601 396 420 14195 14608 25 26 14490 SDFFNSRXL $T=1401620 1303390 0 180 $X=1389660 $Y=1299450
X1844 14150 14582 14659 396 420 13924 14621 25 26 14553 SDFFNSRXL $T=1401620 1325530 0 180 $X=1389660 $Y=1321590
X1845 13942 14615 14645 13998 455 14544 14592 25 26 14742 SDFFNSRXL $T=1390580 1200070 1 0 $X=1390578 $Y=1196130
X1846 13942 14634 14640 13998 14673 14731 14706 25 26 14745 SDFFNSRXL $T=1390580 1214830 0 0 $X=1390578 $Y=1214578
X1847 428 14613 14641 396 459 13890 14660 25 26 465 SDFFNSRXL $T=1390580 1347670 1 0 $X=1390578 $Y=1343730
X1848 14518 14734 14729 13998 418 13671 14633 25 26 14628 SDFFNSRXL $T=1402540 1133650 1 180 $X=1390580 $Y=1133398
X1849 14518 14735 14730 13998 14673 14270 14637 25 26 14611 SDFFNSRXL $T=1402540 1141030 1 180 $X=1390580 $Y=1140778
X1850 14465 14697 14711 13687 438 14496 14635 25 26 14464 SDFFNSRXL $T=1402540 1236970 0 180 $X=1390580 $Y=1233030
X1851 14518 14675 14738 13998 14673 14663 14643 25 26 14622 SDFFNSRXL $T=1403460 1163170 0 180 $X=1391500 $Y=1159230
X1852 14150 14608 14747 396 420 14671 14668 25 26 14550 SDFFNSRXL $T=1404380 1310770 0 180 $X=1392420 $Y=1306830
X1853 14150 14646 14684 396 14673 14149 14778 25 26 14716 SDFFNSRXL $T=1395180 1288630 1 0 $X=1395178 $Y=1284690
X1854 14518 14637 14772 13998 14673 14022 14675 25 26 14672 SDFFNSRXL $T=1407140 1148410 0 180 $X=1395180 $Y=1144470
X1855 14599 14668 14665 396 455 14233 14620 25 26 14840 SDFFNSRXL $T=1397020 1310770 0 0 $X=1397018 $Y=1310518
X1856 14518 14786 14708 13998 14596 13374 14682 25 26 14688 SDFFNSRXL $T=1408980 1170550 1 180 $X=1397020 $Y=1170298
X1857 14465 14777 14771 13687 14596 14405 14697 25 26 14689 SDFFNSRXL $T=1408980 1244350 0 180 $X=1397020 $Y=1240410
X1858 13942 14696 14709 13998 14596 13892 14809 25 26 14788 SDFFNSRXL $T=1398860 1200070 0 0 $X=1398858 $Y=1199818
X1859 14518 14428 14627 13998 455 13690 14612 25 26 14807 SDFFNSRXL $T=1399780 1185310 0 0 $X=1399778 $Y=1185058
X1860 14607 14739 14712 13687 14596 13441 14713 25 26 14813 SDFFNSRXL $T=1400700 1281250 1 0 $X=1400698 $Y=1277310
X1861 14465 14733 14746 13687 14596 14580 14739 25 26 14842 SDFFNSRXL $T=1401160 1259110 0 0 $X=1401158 $Y=1258858
X1862 14599 14782 14846 14810 14673 14546 14754 25 26 14704 SDFFNSRXL $T=1414960 1325530 1 180 $X=1403000 $Y=1325278
X1863 14751 14755 14759 13998 467 14731 14634 25 26 14989 SDFFNSRXL $T=1403460 1214830 0 0 $X=1403458 $Y=1214578
X1864 14599 14760 14775 396 14673 14233 14853 25 26 14818 SDFFNSRXL $T=1403920 1318150 1 0 $X=1403918 $Y=1314210
X1865 14751 14809 14852 13998 469 13738 14755 25 26 14692 SDFFNSRXL $T=1415880 1207450 1 180 $X=1403920 $Y=1207198
X1866 14518 14766 14767 13998 14596 14136 14734 25 26 14843 SDFFNSRXL $T=1404380 1133650 1 0 $X=1404378 $Y=1129710
X1867 14400 14858 14779 14831 406 14403 14761 25 26 14642 SDFFNSRXL $T=1416340 1111510 1 180 $X=1404380 $Y=1111258
X1868 14400 14860 14855 14831 14673 13734 14762 25 26 14756 SDFFNSRXL $T=1416340 1126270 0 180 $X=1404380 $Y=1122330
X1869 14518 14643 14854 14831 14596 13694 14768 25 26 14714 SDFFNSRXL $T=1416340 1155790 0 180 $X=1404380 $Y=1151850
X1870 14837 14844 14856 13998 14673 14544 14770 25 26 14758 SDFFNSRXL $T=1416340 1200070 0 180 $X=1404380 $Y=1196130
X1871 14465 14864 14815 14810 14673 13948 14777 25 26 14764 SDFFNSRXL $T=1416800 1251730 0 180 $X=1404840 $Y=1247790
X1872 14599 14754 14863 14810 14673 13924 14760 25 26 14693 SDFFNSRXL $T=1416800 1318150 1 180 $X=1404840 $Y=1317898
X1873 14599 14578 14861 396 14673 14391 14782 25 26 14776 SDFFNSRXL $T=1418180 1332910 0 180 $X=1406220 $Y=1328970
X1874 14400 14761 14859 14831 469 13906 14766 25 26 14604 SDFFNSRXL $T=1418640 1118890 1 180 $X=1406680 $Y=1118638
X1875 14518 14762 14799 14831 14596 13671 14735 25 26 14890 SDFFNSRXL $T=1407600 1133650 0 0 $X=1407598 $Y=1133398
X1876 14518 14796 14769 13998 14596 13690 14781 25 26 14800 SDFFNSRXL $T=1407600 1185310 1 0 $X=1407598 $Y=1181370
X1877 14868 14797 14877 14831 14596 14663 14795 25 26 14787 SDFFNSRXL $T=1419560 1163170 0 180 $X=1407600 $Y=1159230
X1878 14607 14802 14880 14810 469 14801 14792 25 26 14690 SDFFNSRXL $T=1419560 1266490 0 180 $X=1407600 $Y=1262550
X1879 14607 14713 14808 14810 14673 14149 14886 25 26 14753 SDFFNSRXL $T=1408060 1288630 1 0 $X=1408058 $Y=1284690
X1880 14607 14885 14882 14810 14673 14801 14802 25 26 14699 SDFFNSRXL $T=1420020 1266490 1 180 $X=1408060 $Y=1266238
X1881 14518 14781 14888 14865 14596 13374 14806 25 26 14783 SDFFNSRXL $T=1420940 1170550 1 180 $X=1408980 $Y=1170298
X1882 14607 14851 14895 14810 14673 14671 14835 25 26 14803 SDFFNSRXL $T=1422320 1303390 1 180 $X=1410360 $Y=1303138
X1883 14518 14806 14841 14831 14596 14839 14786 25 26 14644 SDFFNSRXL $T=1422780 1170550 0 180 $X=1410820 $Y=1166610
X1884 14607 14886 14899 14810 469 13736 14834 25 26 14784 SDFFNSRXL $T=1422780 1296010 0 180 $X=1410820 $Y=1292070
X1885 14607 14835 14912 14810 469 14502 14636 25 26 14678 SDFFNSRXL $T=1423240 1296010 1 180 $X=1411280 $Y=1295758
X1886 14751 14792 14850 14810 14596 13660 14920 25 26 14884 SDFFNSRXL $T=1412200 1251730 0 0 $X=1412198 $Y=1251478
X1887 14868 14914 14832 14865 14673 13354 14796 25 26 14774 SDFFNSRXL $T=1424620 1177930 1 180 $X=1412660 $Y=1177678
X1888 14837 14889 14866 14865 14673 13892 14844 25 26 14702 SDFFNSRXL $T=1424620 1200070 1 180 $X=1412660 $Y=1199818
X1889 14751 14862 14873 14865 14596 14496 14849 25 26 14812 SDFFNSRXL $T=1424620 1229590 1 180 $X=1412660 $Y=1229338
X1890 14751 14920 14916 14810 14596 14405 14862 25 26 14848 SDFFNSRXL $T=1426460 1244350 0 180 $X=1414500 $Y=1240410
X1891 14868 14795 14878 14831 478 13735 14950 25 26 14974 SDFFNSRXL $T=1416340 1163170 0 0 $X=1416338 $Y=1162918
X1892 14868 14981 14951 14865 478 14544 14889 25 26 14883 SDFFNSRXL $T=1430140 1200070 0 180 $X=1418180 $Y=1196130
X1893 14599 14941 14900 483 14673 13391 476 25 26 14785 SDFFNSRXL $T=1431060 1340290 0 180 $X=1419100 $Y=1336350
X1894 14751 14817 14915 14865 482 13738 14939 25 26 14988 SDFFNSRXL $T=1420020 1214830 1 0 $X=1420018 $Y=1210890
X1895 14284 14949 14943 14831 469 13677 14858 25 26 14893 SDFFNSRXL $T=1432440 1118890 0 180 $X=1420480 $Y=1114950
X1896 14607 14881 14959 14810 14596 13441 14898 25 26 14871 SDFFNSRXL $T=1432440 1281250 0 180 $X=1420480 $Y=1277310
X1897 14868 14919 14925 14831 482 14663 14928 25 26 15017 SDFFNSRXL $T=1420940 1155790 0 0 $X=1420938 $Y=1155538
X1898 14868 14994 14990 14865 469 13374 14914 25 26 14752 SDFFNSRXL $T=1432900 1170550 1 180 $X=1420940 $Y=1170298
X1899 14518 14922 14927 14831 14673 14270 15012 25 26 14924 SDFFNSRXL $T=1421400 1141030 0 0 $X=1421398 $Y=1140778
X1900 14751 15013 14991 14865 469 13744 14923 25 26 14763 SDFFNSRXL $T=1433360 1229590 0 180 $X=1421400 $Y=1225650
X1901 14868 14816 14931 14865 486 14623 14957 25 26 15117 SDFFNSRXL $T=1421860 1192690 1 0 $X=1421858 $Y=1188750
X1902 14751 14930 14933 14810 467 13746 15019 25 26 15021 SDFFNSRXL $T=1422320 1244350 0 0 $X=1422318 $Y=1244098
X1903 14751 14923 14972 14865 469 14496 14930 25 26 14791 SDFFNSRXL $T=1434740 1236970 0 180 $X=1422780 $Y=1233030
X1904 14599 15023 14982 14810 467 13924 14938 25 26 14934 SDFFNSRXL $T=1435660 1325530 0 180 $X=1423700 $Y=1321590
X1905 14751 14945 14891 14810 478 13660 14864 25 26 15048 SDFFNSRXL $T=1424160 1251730 0 0 $X=1424158 $Y=1251478
X1906 14284 15012 14986 14831 469 14136 14944 25 26 14811 SDFFNSRXL $T=1436120 1133650 0 180 $X=1424160 $Y=1129710
X1907 14751 15019 15026 14810 469 14580 14946 25 26 14845 SDFFNSRXL $T=1436120 1259110 0 180 $X=1424160 $Y=1255170
X1908 14751 14946 14947 14810 469 13707 14885 25 26 14857 SDFFNSRXL $T=1436120 1259110 1 180 $X=1424160 $Y=1258858
X1909 14599 15027 14997 483 469 14391 14941 25 26 14798 SDFFNSRXL $T=1436120 1332910 1 180 $X=1424160 $Y=1332658
X1910 14868 14950 14956 14831 467 14839 14994 25 26 15039 SDFFNSRXL $T=1424620 1170550 1 0 $X=1424618 $Y=1166610
X1911 14607 14952 14948 14810 467 13736 15031 25 26 15072 SDFFNSRXL $T=1424620 1296010 1 0 $X=1424618 $Y=1292070
X1912 14599 14953 14960 14810 487 14233 15014 25 26 15070 SDFFNSRXL $T=1424620 1310770 0 0 $X=1424618 $Y=1310518
X1913 14284 15030 15024 14831 469 14403 14949 25 26 14687 SDFFNSRXL $T=1436580 1111510 1 180 $X=1424620 $Y=1111258
X1914 14284 14944 14935 14831 469 13734 14860 25 26 14597 SDFFNSRXL $T=1436580 1126270 1 180 $X=1424620 $Y=1126018
X1915 14607 15014 14984 14810 467 14671 14945 25 26 14940 SDFFNSRXL $T=1436580 1303390 1 180 $X=1424620 $Y=1303138
X1916 14868 14954 14967 14865 486 13354 15034 25 26 15071 SDFFNSRXL $T=1425080 1177930 0 0 $X=1425078 $Y=1177678
X1917 14868 14957 14963 14865 467 13690 14954 25 26 15037 SDFFNSRXL $T=1425080 1185310 1 0 $X=1425078 $Y=1181370
X1918 14751 14958 14964 14865 478 13875 15013 25 26 15077 SDFFNSRXL $T=1425080 1222210 1 0 $X=1425078 $Y=1218270
X1919 14599 14938 14965 14810 478 13741 15027 25 26 15073 SDFFNSRXL $T=1425080 1325530 0 0 $X=1425078 $Y=1325278
X1920 14599 14969 14971 483 467 15035 15041 25 26 15166 SDFFNSRXL $T=1426000 1340290 0 0 $X=1425998 $Y=1340038
X1921 14284 14976 14979 14831 482 14022 14922 25 26 15063 SDFFNSRXL $T=1427380 1148410 1 0 $X=1427378 $Y=1144470
X1922 14284 14928 14980 14831 478 14022 14976 25 26 15076 SDFFNSRXL $T=1427380 1148410 0 0 $X=1427378 $Y=1148158
X1923 484 14977 14983 483 467 13890 14969 25 26 15061 SDFFNSRXL $T=1427380 1347670 1 0 $X=1427378 $Y=1343730
X1924 14751 14939 14987 14865 467 13738 14981 25 26 14995 SDFFNSRXL $T=1428300 1207450 0 0 $X=1428298 $Y=1207198
X1925 14868 15058 15055 14831 491 13735 14919 25 26 14978 SDFFNSRXL $T=1440260 1163170 1 180 $X=1428300 $Y=1162918
X1926 14607 15068 14996 14810 478 14581 14952 25 26 14985 SDFFNSRXL $T=1441180 1281250 1 180 $X=1429220 $Y=1280998
X1927 15135 15123 15042 14865 482 14838 14958 25 26 15018 SDFFNSRXL $T=1444860 1222210 1 180 $X=1432900 $Y=1221958
X1928 14751 15113 15052 14810 482 13746 15032 25 26 15025 SDFFNSRXL $T=1446240 1244350 1 180 $X=1434280 $Y=1244098
X1929 494 15147 15074 483 478 444 14977 25 26 15033 SDFFNSRXL $T=1447620 1347670 1 180 $X=1435660 $Y=1347418
X1930 14607 15040 15060 14810 482 13441 15086 25 26 15067 SDFFNSRXL $T=1437500 1281250 1 0 $X=1437498 $Y=1277310
X1931 14868 15129 15064 14865 491 13712 15056 25 26 14975 SDFFNSRXL $T=1449920 1192690 1 180 $X=1437960 $Y=1192438
X1932 14284 15115 15167 14831 499 14403 15062 25 26 15054 SDFFNSRXL $T=1450380 1111510 1 180 $X=1438420 $Y=1111258
X1933 14751 15078 15084 14865 500 13745 15083 25 26 15119 SDFFNSRXL $T=1439800 1236970 0 0 $X=1439798 $Y=1236718
X1934 14284 15201 15122 14831 488 14136 14962 25 26 15069 SDFFNSRXL $T=1451760 1133650 0 180 $X=1439800 $Y=1129710
X1935 14284 15062 15165 14831 491 14022 15080 25 26 15046 SDFFNSRXL $T=1452220 1148410 0 180 $X=1440260 $Y=1144470
X1936 14868 15034 15091 14865 486 13354 15058 25 26 15235 SDFFNSRXL $T=1440720 1177930 0 0 $X=1440718 $Y=1177678
X1937 14751 15032 15107 14810 488 14405 15078 25 26 15163 SDFFNSRXL $T=1440720 1244350 1 0 $X=1440718 $Y=1240410
X1938 14284 15090 15111 14831 499 13671 15201 25 26 15160 SDFFNSRXL $T=1441180 1133650 0 0 $X=1441178 $Y=1133398
X1939 14284 15080 15112 14831 482 14022 15090 25 26 15240 SDFFNSRXL $T=1441180 1148410 0 0 $X=1441178 $Y=1148158
X1940 14607 15086 15114 14810 500 14581 15068 25 26 15219 SDFFNSRXL $T=1441180 1281250 0 0 $X=1441178 $Y=1280998
X1941 14607 15031 15087 14810 487 14502 15081 25 26 15049 SDFFNSRXL $T=1441640 1296010 0 0 $X=1441638 $Y=1295758
X1942 15135 15210 15164 14810 491 13707 15113 25 26 15043 SDFFNSRXL $T=1453600 1259110 1 180 $X=1441640 $Y=1258858
X1943 14599 504 15124 14810 478 14233 14953 25 26 15089 SDFFNSRXL $T=1453600 1318150 0 180 $X=1441640 $Y=1314210
X1944 14284 15214 15200 14831 503 13906 15115 25 26 15106 SDFFNSRXL $T=1454060 1118890 1 180 $X=1442100 $Y=1118638
X1945 15225 15081 15212 14810 482 14195 15118 25 26 15088 SDFFNSRXL $T=1454060 1303390 0 180 $X=1442100 $Y=1299450
X1946 14868 15226 15116 14865 488 13712 15129 25 26 15127 SDFFNSRXL $T=1455440 1192690 0 180 $X=1443480 $Y=1188750
X1947 15135 15056 15092 14865 491 13738 15120 25 26 15047 SDFFNSRXL $T=1455440 1207450 1 180 $X=1443480 $Y=1207198
X1948 15135 15120 15146 14865 488 14838 15123 25 26 15252 SDFFNSRXL $T=1444860 1222210 0 0 $X=1444858 $Y=1221958
X1949 14868 15145 15153 14865 486 14623 15226 25 26 15261 SDFFNSRXL $T=1445320 1185310 0 0 $X=1445318 $Y=1185058
X1950 15135 15258 15222 14810 499 13746 15154 25 26 15150 SDFFNSRXL $T=1458200 1244350 1 180 $X=1446240 $Y=1244098
X1951 15135 15083 15199 14865 500 14496 15248 25 26 15268 SDFFNSRXL $T=1448540 1229590 0 0 $X=1448538 $Y=1229338
X1952 15225 15108 15286 14810 482 13741 15197 25 26 15157 SDFFNSRXL $T=1460960 1325530 1 180 $X=1449000 $Y=1325278
X1953 15135 15242 15237 14810 486 14801 15210 25 26 15355 SDFFNSRXL $T=1454520 1266490 1 0 $X=1454518 $Y=1262550
X1954 494 15243 15245 483 500 15035 505 25 26 15344 SDFFNSRXL $T=1454520 1340290 1 0 $X=1454518 $Y=1336350
X1955 15353 15260 15346 14831 511 13734 15214 25 26 15159 SDFFNSRXL $T=1466480 1126270 0 180 $X=1454520 $Y=1122330
X1956 15358 15267 15345 14831 15321 13735 15238 25 26 15161 SDFFNSRXL $T=1466480 1163170 1 180 $X=1454520 $Y=1162918
X1957 15135 15249 15257 14810 486 13534 15314 25 26 15361 SDFFNSRXL $T=1454980 1273870 1 0 $X=1454978 $Y=1269930
X1958 15358 15272 15294 14831 15321 13735 15244 25 26 15202 SDFFNSRXL $T=1466940 1163170 0 180 $X=1454980 $Y=1159230
X1959 15225 15350 15349 14810 512 14671 15254 25 26 15221 SDFFNSRXL $T=1466940 1303390 1 180 $X=1454980 $Y=1303138
X1960 15135 15255 15263 14865 15321 13738 15262 25 26 15287 SDFFNSRXL $T=1455440 1207450 0 0 $X=1455438 $Y=1207198
X1961 15353 15278 15343 14831 511 14136 15260 25 26 15139 SDFFNSRXL $T=1468320 1133650 0 180 $X=1456360 $Y=1129710
X1962 15135 15248 15279 14865 499 13745 15370 25 26 15288 SDFFNSRXL $T=1456820 1236970 1 0 $X=1456818 $Y=1233030
X1963 15135 15154 15276 14810 503 13660 15371 25 26 15218 SDFFNSRXL $T=1456820 1251730 0 0 $X=1456818 $Y=1251478
X1964 14868 15324 15270 14865 503 13892 15273 25 26 15066 SDFFNSRXL $T=1468780 1200070 1 180 $X=1456820 $Y=1199818
X1965 14284 15274 15283 14831 478 13694 15272 25 26 15356 SDFFNSRXL $T=1457280 1155790 1 0 $X=1457278 $Y=1151850
X1966 15353 15368 15364 14831 503 13671 15278 25 26 15192 SDFFNSRXL $T=1469240 1133650 1 180 $X=1457280 $Y=1133398
X1967 15358 15295 15275 14865 15321 14586 15267 25 26 15216 SDFFNSRXL $T=1469240 1177930 0 180 $X=1457280 $Y=1173990
X1968 15358 15316 15365 14865 499 14623 15145 25 26 15082 SDFFNSRXL $T=1469240 1185310 1 180 $X=1457280 $Y=1185058
X1969 15292 15369 15277 15340 488 14466 15249 25 26 15266 SDFFNSRXL $T=1469240 1273870 1 180 $X=1457280 $Y=1273618
X1970 15135 15379 15366 15340 500 13948 15258 25 26 15170 SDFFNSRXL $T=1470160 1244350 1 180 $X=1458200 $Y=1244098
X1971 15292 15254 15351 15340 499 14195 15285 25 26 15281 SDFFNSRXL $T=1470160 1303390 0 180 $X=1458200 $Y=1299450
X1972 14284 15291 15312 14831 511 13906 15368 25 26 15409 SDFFNSRXL $T=1458660 1118890 0 0 $X=1458658 $Y=1118638
X1973 15135 15370 15378 14865 503 14838 15289 25 26 15284 SDFFNSRXL $T=1470620 1222210 1 180 $X=1458660 $Y=1221958
X1974 14599 15197 15362 483 482 14391 15298 25 26 15151 SDFFNSRXL $T=1470620 1332910 1 180 $X=1458660 $Y=1332658
X1975 15358 15384 15382 14865 515 13690 15295 25 26 15234 SDFFNSRXL $T=1471080 1185310 0 180 $X=1459120 $Y=1181370
X1976 15293 15320 15323 14831 499 14403 15291 25 26 15407 SDFFNSRXL $T=1459580 1111510 0 0 $X=1459578 $Y=1111258
X1977 15353 15399 15337 14831 516 14270 15274 25 26 15168 SDFFNSRXL $T=1471540 1141030 1 180 $X=1459580 $Y=1140778
X1978 15358 15244 15359 14865 15321 13374 15316 25 26 15194 SDFFNSRXL $T=1471540 1170550 1 180 $X=1459580 $Y=1170298
X1979 15353 15262 15401 14865 15321 14691 15324 25 26 15317 SDFFNSRXL $T=1472000 1207450 0 180 $X=1460040 $Y=1203510
X1980 494 522 15381 483 488 444 15147 25 26 15319 SDFFNSRXL $T=1472000 1347670 1 180 $X=1460040 $Y=1347418
X1981 15437 15314 15380 15340 519 14801 15242 25 26 15280 SDFFNSRXL $T=1472460 1266490 1 180 $X=1460500 $Y=1266238
X1982 15292 15285 15332 15340 15321 14581 15369 25 26 15363 SDFFNSRXL $T=1460960 1281250 0 0 $X=1460958 $Y=1280998
X1983 14868 15273 15338 14865 15321 13712 15373 25 26 15375 SDFFNSRXL $T=1461880 1192690 0 0 $X=1461878 $Y=1192438
X1984 15225 15118 15412 14810 488 14671 15334 25 26 15282 SDFFNSRXL $T=1473840 1310770 0 180 $X=1461880 $Y=1306830
X1985 15225 15334 15341 14810 499 14233 15036 25 26 15239 SDFFNSRXL $T=1473840 1310770 1 180 $X=1461880 $Y=1310518
X1986 15225 15298 15342 14810 519 13741 15416 25 26 15442 SDFFNSRXL $T=1462800 1325530 0 0 $X=1462798 $Y=1325278
X1987 15292 15479 15415 15340 503 14502 15350 25 26 15377 SDFFNSRXL $T=1480280 1296010 1 180 $X=1468320 $Y=1295758
X1988 15293 15398 15403 14831 488 13671 15399 25 26 15503 SDFFNSRXL $T=1469240 1133650 0 0 $X=1469238 $Y=1133398
X1989 15293 15424 15446 14831 491 14022 15405 25 26 15325 SDFFNSRXL $T=1482120 1148410 0 180 $X=1470160 $Y=1144470
X1990 15225 15509 15507 14810 500 13924 15406 25 26 15265 SDFFNSRXL $T=1482580 1318150 0 180 $X=1470620 $Y=1314210
X1991 15358 15420 15425 14865 478 14586 15486 25 26 15528 SDFFNSRXL $T=1472000 1170550 0 0 $X=1471998 $Y=1170298
X1992 15353 15421 15426 14865 486 13744 15455 25 26 15526 SDFFNSRXL $T=1472000 1229590 1 0 $X=1471998 $Y=1225650
X1993 15358 15373 15431 14865 478 14623 15420 25 26 15521 SDFFNSRXL $T=1472460 1185310 0 0 $X=1472458 $Y=1185058
X1994 15292 15423 15429 15340 482 14466 15449 25 26 15456 SDFFNSRXL $T=1472460 1273870 0 0 $X=1472458 $Y=1273618
X1995 15293 15428 15438 14831 503 14403 15320 25 26 15537 SDFFNSRXL $T=1472920 1111510 1 0 $X=1472918 $Y=1107570
X1996 15292 14778 15441 15340 512 14149 15524 25 26 15339 SDFFNSRXL $T=1472920 1288630 1 0 $X=1472918 $Y=1284690
X1997 15358 15508 15430 14831 515 14839 15424 25 26 15228 SDFFNSRXL $T=1484880 1163170 1 180 $X=1472920 $Y=1162918
X1998 15292 15524 15457 15340 519 13736 15243 25 26 15376 SDFFNSRXL $T=1484880 1296010 0 180 $X=1472920 $Y=1292070
X1999 494 15525 15445 483 512 15035 15434 25 26 15372 SDFFNSRXL $T=1484880 1340290 1 180 $X=1472920 $Y=1340038
X2000 15353 15329 15443 14865 482 13875 15421 25 26 15551 SDFFNSRXL $T=1473380 1222210 1 0 $X=1473378 $Y=1218270
X2001 15225 15406 15452 14810 488 14671 15538 25 26 15609 SDFFNSRXL $T=1473840 1310770 1 0 $X=1473838 $Y=1306830
X2002 494 15472 528 483 512 444 525 25 26 524 SDFFNSRXL $T=1485800 1347670 1 180 $X=1473840 $Y=1347418
X2003 15135 15440 15459 15340 527 13660 15541 25 26 15488 SDFFNSRXL $T=1474760 1251730 0 0 $X=1474758 $Y=1251478
X2004 15225 15416 15461 14810 15321 13741 15477 25 26 15433 SDFFNSRXL $T=1474760 1325530 0 0 $X=1474758 $Y=1325278
X2005 15292 15541 15460 15340 15321 13534 15423 25 26 15264 SDFFNSRXL $T=1486720 1266490 1 180 $X=1474760 $Y=1266238
X2006 14868 15458 15465 14865 482 13712 15400 25 26 15545 SDFFNSRXL $T=1475220 1192690 0 0 $X=1475218 $Y=1192438
X2007 15225 15434 15467 483 488 15035 15485 25 26 15611 SDFFNSRXL $T=1475220 1340290 1 0 $X=1475218 $Y=1336350
X2008 15353 15405 15436 14831 482 14270 15413 25 26 15504 SDFFNSRXL $T=1476600 1141030 0 0 $X=1476598 $Y=1140778
X2009 15292 15449 15473 15340 527 13534 15556 25 26 15483 SDFFNSRXL $T=1476600 1273870 1 0 $X=1476598 $Y=1269930
X2010 15293 15453 15530 14831 499 13906 15468 25 26 15464 SDFFNSRXL $T=1488560 1118890 1 180 $X=1476600 $Y=1118638
X2011 15353 15549 15540 14865 515 14544 15458 25 26 15360 SDFFNSRXL $T=1488560 1200070 0 180 $X=1476600 $Y=1196130
X2012 15353 15550 15529 14865 516 14691 15471 25 26 15357 SDFFNSRXL $T=1488560 1207450 0 180 $X=1476600 $Y=1203510
X2013 15437 15335 15422 15340 482 14580 15440 25 26 15466 SDFFNSRXL $T=1488560 1259110 0 180 $X=1476600 $Y=1255170
X2014 494 15485 15546 483 499 13890 15472 25 26 15354 SDFFNSRXL $T=1488560 1347670 0 180 $X=1476600 $Y=1343730
X2015 15293 15474 15475 14831 511 13734 15398 25 26 15612 SDFFNSRXL $T=1477520 1126270 0 0 $X=1477518 $Y=1126018
X2016 15358 15486 15490 14831 478 13735 15557 25 26 15531 SDFFNSRXL $T=1478900 1163170 1 0 $X=1478898 $Y=1159230
X2017 15358 15238 15543 14831 516 14839 15508 25 26 15203 SDFFNSRXL $T=1492240 1170550 0 180 $X=1480280 $Y=1166610
X2018 15225 15538 15542 15340 515 14502 15506 25 26 15411 SDFFNSRXL $T=1492240 1296010 1 180 $X=1480280 $Y=1295758
X2019 14732 15512 15518 14865 499 14731 15550 25 26 15670 SDFFNSRXL $T=1480740 1214830 1 0 $X=1480738 $Y=1210890
X2020 15225 15489 15533 14810 500 13924 15509 25 26 15625 SDFFNSRXL $T=1482580 1318150 1 0 $X=1482578 $Y=1314210
X2021 15293 15468 15536 14831 499 14403 15428 25 26 15635 SDFFNSRXL $T=1483040 1111510 0 0 $X=1483038 $Y=1111258
X2022 15358 15557 15561 14831 491 14663 15627 25 26 15482 SDFFNSRXL $T=1487180 1155790 0 0 $X=1487178 $Y=1155538
X2023 14732 15671 15575 15340 491 14838 15512 25 26 15555 SDFFNSRXL $T=1499600 1222210 0 180 $X=1487640 $Y=1218270
X2024 15353 15642 15567 14865 491 14544 15549 25 26 15558 SDFFNSRXL $T=1500980 1192690 1 180 $X=1489020 $Y=1192438
X2025 494 532 15577 534 499 13890 15696 25 26 15652 SDFFNSRXL $T=1489480 1347670 1 0 $X=1489478 $Y=1343730
X2026 15293 15570 15595 14831 499 13906 15616 25 26 15669 SDFFNSRXL $T=1489940 1118890 0 0 $X=1489938 $Y=1118638
X2027 15292 15572 15599 15340 491 14149 15617 25 26 15432 SDFFNSRXL $T=1489940 1288630 0 0 $X=1489938 $Y=1288378
X2028 15293 15627 15646 14831 491 14270 15574 25 26 15480 SDFFNSRXL $T=1502360 1141030 1 180 $X=1490400 $Y=1140778
X2029 15358 15600 15610 14865 15321 14586 15640 25 26 15757 SDFFNSRXL $T=1490860 1170550 0 0 $X=1490858 $Y=1170298
X2030 14732 15719 15711 14865 515 14691 15601 25 26 15447 SDFFNSRXL $T=1502820 1207450 0 180 $X=1490860 $Y=1203510
X2031 15760 15720 15596 15340 491 14580 15602 25 26 15444 SDFFNSRXL $T=1502820 1259110 0 180 $X=1490860 $Y=1255170
X2032 15292 15607 15613 15340 512 14466 15572 25 26 15742 SDFFNSRXL $T=1491320 1273870 0 0 $X=1491318 $Y=1273618
X2033 15631 15694 15634 15340 527 13948 15604 25 26 15597 SDFFNSRXL $T=1503280 1244350 1 180 $X=1491320 $Y=1244098
X2034 15293 15616 15620 14831 503 13734 15474 25 26 15562 SDFFNSRXL $T=1503740 1126270 0 180 $X=1491780 $Y=1122330
X2035 544 542 541 534 499 444 532 25 26 531 SDFFNSRXL $T=1503740 1347670 1 180 $X=1491780 $Y=1347418
X2036 15437 15514 15565 15340 527 13745 15462 25 26 15630 SDFFNSRXL $T=1492240 1236970 1 0 $X=1492238 $Y=1233030
X2037 15225 15619 15618 534 503 13741 15632 25 26 15668 SDFFNSRXL $T=1492240 1325530 0 0 $X=1492238 $Y=1325278
X2038 15292 15737 15608 15340 15321 13736 15479 25 26 15402 SDFFNSRXL $T=1504660 1296010 0 180 $X=1492700 $Y=1292070
X2039 15437 15602 15638 15340 503 14580 15694 25 26 15756 SDFFNSRXL $T=1493160 1251730 0 0 $X=1493158 $Y=1251478
X2040 15358 15574 15647 14831 515 13735 15600 25 26 15751 SDFFNSRXL $T=1494080 1163170 1 0 $X=1494078 $Y=1159230
X2041 15631 15639 15649 15340 538 13707 15720 25 26 15717 SDFFNSRXL $T=1494080 1259110 0 0 $X=1494078 $Y=1258858
X2042 15292 15556 15650 15340 503 14466 15607 25 26 15754 SDFFNSRXL $T=1494080 1273870 1 0 $X=1494078 $Y=1269930
X2043 15293 15745 15690 14831 503 13677 15570 25 26 15628 SDFFNSRXL $T=1506040 1118890 0 180 $X=1494080 $Y=1114950
X2044 15353 15601 15733 15687 503 13892 15637 25 26 15629 SDFFNSRXL $T=1506040 1200070 1 180 $X=1494080 $Y=1199818
X2045 15225 15746 15712 534 15321 13924 15645 25 26 15469 SDFFNSRXL $T=1506040 1318150 1 180 $X=1494080 $Y=1317898
X2046 544 15696 15621 534 500 15035 15525 25 26 15626 SDFFNSRXL $T=1506040 1340290 1 180 $X=1494080 $Y=1340038
X2047 15292 15662 15681 15340 519 14195 15737 25 26 15740 SDFFNSRXL $T=1497760 1303390 1 0 $X=1497758 $Y=1299450
X2048 15760 15605 15854 15340 538 14581 15749 25 26 15689 SDFFNSRXL $T=1516160 1281250 0 180 $X=1504200 $Y=1277310
X2049 15631 15774 15779 15340 503 14405 15848 25 26 15803 SDFFNSRXL $T=1506500 1236970 1 0 $X=1506498 $Y=1233030
X2050 15631 15604 15783 15340 548 13948 15774 25 26 15880 SDFFNSRXL $T=1506960 1244350 0 0 $X=1506958 $Y=1244098
X2051 15358 15762 15786 15687 15321 14586 15857 25 26 15734 SDFFNSRXL $T=1507420 1177930 1 0 $X=1507418 $Y=1173990
X2052 15926 15873 15785 15687 515 14839 15762 25 26 15775 SDFFNSRXL $T=1519380 1170550 0 180 $X=1507420 $Y=1166610
X2053 544 15796 15794 534 15321 13924 15746 25 26 15755 SDFFNSRXL $T=1519380 1318150 0 180 $X=1507420 $Y=1314210
X2054 544 15841 15870 534 515 15035 15782 25 26 15766 SDFFNSRXL $T=1519380 1340290 0 180 $X=1507420 $Y=1336350
X2055 544 15829 552 534 549 547 545 25 26 543 SDFFNSRXL $T=1519380 1347670 1 180 $X=1507420 $Y=1347418
X2056 14732 15840 15788 15687 511 14731 15671 25 26 15688 SDFFNSRXL $T=1519840 1214830 0 180 $X=1507880 $Y=1210890
X2057 15293 15793 15797 15687 516 14022 15853 25 26 15867 SDFFNSRXL $T=1508340 1141030 0 0 $X=1508338 $Y=1140778
X2058 14732 15834 15787 15687 538 14731 15795 25 26 15723 SDFFNSRXL $T=1520300 1207450 1 180 $X=1508340 $Y=1207198
X2059 544 15828 15878 534 15321 14671 15796 25 26 15727 SDFFNSRXL $T=1520760 1310770 0 180 $X=1508800 $Y=1306830
X2060 15292 15813 15798 15340 511 14502 15849 25 26 15724 SDFFNSRXL $T=1510180 1288630 0 0 $X=1510178 $Y=1288378
X2061 15760 15827 15843 15340 548 14801 15901 25 26 15860 SDFFNSRXL $T=1510640 1259110 0 0 $X=1510638 $Y=1258858
X2062 15926 15835 15801 15687 511 14136 15808 25 26 15682 SDFFNSRXL $T=1522600 1126270 1 180 $X=1510640 $Y=1126018
X2063 15926 15896 15876 15687 516 14663 15793 25 26 15715 SDFFNSRXL $T=1522600 1148410 1 180 $X=1510640 $Y=1148158
X2064 15937 15857 15890 15687 516 14623 15833 25 26 15790 SDFFNSRXL $T=1522600 1185310 0 180 $X=1510640 $Y=1181370
X2065 14732 15856 15877 15687 515 13892 15834 25 26 15753 SDFFNSRXL $T=1522600 1200070 0 180 $X=1510640 $Y=1196130
X2066 544 15849 15891 15340 515 14195 15828 25 26 15773 SDFFNSRXL $T=1522600 1303390 0 180 $X=1510640 $Y=1299450
X2067 544 15782 15886 534 549 15035 15829 25 26 15695 SDFFNSRXL $T=1522600 1340290 1 180 $X=1510640 $Y=1340038
X2068 15358 15767 15844 15687 15321 14839 15896 25 26 15836 SDFFNSRXL $T=1511100 1163170 1 0 $X=1511098 $Y=1159230
X2069 15926 15777 15898 15687 538 14136 15835 25 26 15713 SDFFNSRXL $T=1523060 1133650 0 180 $X=1511100 $Y=1129710
X2070 14732 15795 15899 15687 538 14691 15839 25 26 15685 SDFFNSRXL $T=1523060 1207450 0 180 $X=1511100 $Y=1203510
X2071 15937 15916 15900 15340 515 13875 15719 25 26 15826 SDFFNSRXL $T=1523060 1214830 1 180 $X=1511100 $Y=1214578
X2072 15631 15901 15812 15340 511 14580 15639 25 26 15732 SDFFNSRXL $T=1523060 1251730 1 180 $X=1511100 $Y=1251478
X2073 544 15632 15902 534 549 14391 15841 25 26 15741 SDFFNSRXL $T=1523060 1332910 0 180 $X=1511100 $Y=1328970
X2074 15293 15808 15846 15687 503 13906 15745 25 26 15770 SDFFNSRXL $T=1511560 1118890 0 0 $X=1511558 $Y=1118638
X2075 14732 15842 15802 15340 511 14838 15840 25 26 15716 SDFFNSRXL $T=1523520 1222210 1 180 $X=1511560 $Y=1221958
X2076 15926 15853 15920 15687 538 14270 15847 25 26 15714 SDFFNSRXL $T=1523980 1141030 0 180 $X=1512020 $Y=1137090
X2077 15937 15833 15929 15687 15692 14544 15856 25 26 15805 SDFFNSRXL $T=1525820 1192690 0 180 $X=1513860 $Y=1188750
X2078 15942 15749 15957 15340 555 14581 15813 25 26 15861 SDFFNSRXL $T=1528120 1281250 0 180 $X=1516160 $Y=1277310
X2079 15942 15967 15970 15340 548 14502 15874 25 26 15869 SDFFNSRXL $T=1529040 1296010 0 180 $X=1517080 $Y=1292070
X2080 15926 15847 15936 15687 477 14270 15872 25 26 16072 SDFFNSRXL $T=1523520 1133650 0 0 $X=1523518 $Y=1133398
X2081 15926 15855 15948 15687 15692 14839 16049 25 26 15784 SDFFNSRXL $T=1524440 1163170 1 0 $X=1524438 $Y=1159230
X2082 544 15943 15946 534 548 14502 15967 25 26 16115 SDFFNSRXL $T=1524440 1296010 0 0 $X=1524438 $Y=1295758
X2083 544 15940 15950 534 548 14233 15943 25 26 16076 SDFFNSRXL $T=1524440 1310770 0 0 $X=1524438 $Y=1310518
X2084 15926 16048 15951 15687 516 14663 15931 25 26 15799 SDFFNSRXL $T=1536400 1148410 1 180 $X=1524440 $Y=1148158
X2085 15926 16049 16009 15687 477 14586 15873 25 26 15933 SDFFNSRXL $T=1536400 1170550 0 180 $X=1524440 $Y=1166610
X2086 15942 15962 16037 15340 516 14466 15897 25 26 15868 SDFFNSRXL $T=1536400 1273870 0 180 $X=1524440 $Y=1269930
X2087 15941 16012 15963 534 477 13924 15940 25 26 15934 SDFFNSRXL $T=1536400 1318150 0 180 $X=1524440 $Y=1314210
X2088 15937 15839 15953 15687 477 14691 16052 25 26 16074 SDFFNSRXL $T=1524900 1200070 0 0 $X=1524898 $Y=1199818
X2089 15941 15947 15958 534 548 14391 16012 25 26 16062 SDFFNSRXL $T=1524900 1325530 0 0 $X=1524898 $Y=1325278
X2090 15942 15874 15966 15340 515 14149 16054 25 26 15938 SDFFNSRXL $T=1525360 1288630 1 0 $X=1525358 $Y=1284690
X2091 14732 15982 16010 16011 15692 14838 15954 25 26 15863 SDFFNSRXL $T=1537320 1222210 0 180 $X=1525360 $Y=1218270
X2092 15942 15976 15972 16011 15692 14801 15962 25 26 15881 SDFFNSRXL $T=1537780 1266490 0 180 $X=1525820 $Y=1262550
X2093 15942 16054 16053 16011 516 14149 15965 25 26 15882 SDFFNSRXL $T=1537780 1281250 1 180 $X=1525820 $Y=1280998
X2094 15631 15964 15975 15340 516 14405 16041 25 26 15864 SDFFNSRXL $T=1526740 1236970 0 0 $X=1526738 $Y=1236718
X2095 14732 15987 15969 16011 15692 14496 15964 25 26 15858 SDFFNSRXL $T=1538700 1229590 1 180 $X=1526740 $Y=1229338
X2096 14732 15954 15979 16011 516 14838 15987 25 26 15875 SDFFNSRXL $T=1527200 1222210 0 0 $X=1527198 $Y=1221958
X2097 15937 16052 15961 15687 15692 14623 15956 25 26 15879 SDFFNSRXL $T=1539160 1185310 1 180 $X=1527200 $Y=1185058
X2098 15631 16041 15999 16011 548 13948 15976 25 26 15887 SDFFNSRXL $T=1539620 1244350 1 180 $X=1527660 $Y=1244098
X2099 15937 15956 16058 15687 15996 14544 15982 25 26 15977 SDFFNSRXL $T=1540080 1192690 1 180 $X=1528120 $Y=1192438
X2100 15926 16102 16097 15687 477 14270 15994 25 26 15981 SDFFNSRXL $T=1540540 1141030 0 180 $X=1528580 $Y=1137090
X2101 15937 16103 16031 15687 477 14731 15916 25 26 15983 SDFFNSRXL $T=1540540 1214830 0 180 $X=1528580 $Y=1210890
X2102 14732 16004 16007 16011 15996 14496 16103 25 26 16177 SDFFNSRXL $T=1529500 1229590 1 0 $X=1529498 $Y=1225650
X2103 15941 16006 15988 534 477 444 16005 25 26 16100 SDFFNSRXL $T=1529960 1340290 0 0 $X=1529958 $Y=1340038
X2104 15941 16186 16182 534 477 14233 15947 25 26 16035 SDFFNSRXL $T=1546060 1310770 0 180 $X=1534100 $Y=1306830
X2105 15926 16230 16227 15687 15692 14839 16098 25 26 16092 SDFFNSRXL $T=1550200 1163170 1 180 $X=1538240 $Y=1162918
X2106 15942 16112 16114 16011 15996 14466 16253 25 26 16208 SDFFNSRXL $T=1538700 1273870 0 0 $X=1538698 $Y=1273618
X2107 562 573 16129 534 548 444 16006 25 26 16290 SDFFNSRXL $T=1541460 1347670 1 0 $X=1541458 $Y=1343730
X2108 15941 16161 16173 534 548 14546 16283 25 26 16289 SDFFNSRXL $T=1541920 1318150 1 0 $X=1541918 $Y=1314210
X2109 15942 16283 16091 16011 477 14149 16112 25 26 16130 SDFFNSRXL $T=1553880 1288630 0 180 $X=1541920 $Y=1284690
X2110 15941 16005 16198 534 584 444 590 25 26 581 SDFFNSRXL $T=1543760 1340290 0 0 $X=1543758 $Y=1340038
X2111 15926 16191 16200 15687 477 14663 16102 25 26 16313 SDFFNSRXL $T=1544220 1148410 1 0 $X=1544218 $Y=1144470
X2112 15926 16098 16305 15687 15996 14663 16191 25 26 16187 SDFFNSRXL $T=1556640 1148410 1 180 $X=1544680 $Y=1148158
X2113 15937 16310 16303 16011 15692 14496 16203 25 26 16188 SDFFNSRXL $T=1556640 1222210 1 180 $X=1544680 $Y=1221958
X2114 15937 16203 16220 16011 15692 14838 16325 25 26 16386 SDFFNSRXL $T=1545600 1222210 1 0 $X=1545598 $Y=1218270
X2115 16334 16318 16207 16011 15996 14405 16004 25 26 16201 SDFFNSRXL $T=1557560 1244350 0 180 $X=1545600 $Y=1240410
X2116 16334 15965 16312 16011 15692 14801 16214 25 26 16185 SDFFNSRXL $T=1557560 1259110 1 180 $X=1545600 $Y=1258858
X2117 15941 16215 16315 534 15996 14391 16206 25 26 16204 SDFFNSRXL $T=1557560 1325530 1 180 $X=1545600 $Y=1325278
X2118 15937 16222 16317 15687 15692 14691 16212 25 26 16199 SDFFNSRXL $T=1558020 1200070 0 180 $X=1546060 $Y=1196130
X2119 15937 16325 16324 15687 15692 14731 16222 25 26 16213 SDFFNSRXL $T=1558480 1207450 1 180 $X=1546520 $Y=1207198
X2120 15942 16223 16328 534 15996 14502 580 25 26 16186 SDFFNSRXL $T=1558480 1296010 0 180 $X=1546520 $Y=1292070
X2121 15941 16204 16329 534 15996 14546 16039 25 26 16161 SDFFNSRXL $T=1558480 1318150 1 180 $X=1546520 $Y=1317898
X2122 15941 16332 16330 534 584 15035 578 25 26 16215 SDFFNSRXL $T=1558480 1332910 1 180 $X=1546520 $Y=1332658
X2123 15942 16343 16339 534 15996 14195 16172 25 26 16223 SDFFNSRXL $T=1559400 1296010 1 180 $X=1547440 $Y=1295758
X2124 15926 16372 16367 15687 15692 14839 16230 25 26 16246 SDFFNSRXL $T=1562160 1163170 1 180 $X=1550200 $Y=1162918
X2125 15942 16253 16279 16011 15996 14581 16387 25 26 16363 SDFFNSRXL $T=1550660 1273870 0 0 $X=1550658 $Y=1273618
X2126 15937 16358 16440 16011 15996 14496 16202 25 26 16310 SDFFNSRXL $T=1568600 1222210 1 180 $X=1556640 $Y=1221958
X2127 16334 16433 16450 16011 15996 14801 16178 25 26 16340 SDFFNSRXL $T=1570440 1259110 1 180 $X=1558480 $Y=1258858
X2128 16334 16362 16370 16011 15692 14801 16433 25 26 16356 SDFFNSRXL $T=1558940 1266490 1 0 $X=1558938 $Y=1262550
X2129 562 582 16371 534 584 547 597 25 26 16396 SDFFNSRXL $T=1558940 1347670 0 0 $X=1558938 $Y=1347418
X2130 15941 16388 16415 534 15996 14546 563 25 26 16349 SDFFNSRXL $T=1570900 1318150 0 180 $X=1558940 $Y=1314210
X2131 15926 16368 16374 15687 15692 14623 16420 25 26 16446 SDFFNSRXL $T=1559400 1185310 1 0 $X=1559398 $Y=1181370
X2132 16334 16364 16425 16011 584 14405 16333 25 26 16358 SDFFNSRXL $T=1571360 1236970 0 180 $X=1559400 $Y=1233030
X2133 16334 16444 16454 16011 15692 14405 16364 25 26 16359 SDFFNSRXL $T=1571360 1244350 0 180 $X=1559400 $Y=1240410
X2134 15937 16468 16406 15687 584 14731 16183 25 26 16369 SDFFNSRXL $T=1572280 1207450 1 180 $X=1560320 $Y=1207198
X2135 15942 16394 16398 534 584 14671 16455 25 26 16343 SDFFNSRXL $T=1561240 1296010 0 0 $X=1561238 $Y=1295758
X2136 15941 16399 16456 595 15996 14546 16344 25 26 16388 SDFFNSRXL $T=1573200 1325530 0 180 $X=1561240 $Y=1321590
X2137 15937 16391 16404 15687 584 14544 16205 25 26 16390 SDFFNSRXL $T=1562620 1192690 0 0 $X=1562618 $Y=1192438
X2138 562 16396 16419 595 584 444 600 25 26 16332 SDFFNSRXL $T=1562620 1340290 0 0 $X=1562618 $Y=1340038
X2139 15937 16369 16405 15687 584 14691 16389 25 26 16391 SDFFNSRXL $T=1574580 1200070 1 180 $X=1562620 $Y=1199818
X2140 15941 16482 16469 595 584 15035 594 25 26 16399 SDFFNSRXL $T=1574580 1332910 1 180 $X=1562620 $Y=1332658
X2141 16334 16413 16422 16011 584 14580 16280 25 26 16412 SDFFNSRXL $T=1563080 1251730 1 0 $X=1563078 $Y=1247790
X2142 15926 16420 16424 15687 15692 14586 16463 25 26 16411 SDFFNSRXL $T=1563540 1177930 1 0 $X=1563538 $Y=1173990
X2143 15937 16212 16430 15687 584 14691 16170 25 26 16509 SDFFNSRXL $T=1564000 1200070 1 0 $X=1563998 $Y=1196130
X2144 15937 16417 16431 15687 15996 14731 16345 25 26 16468 SDFFNSRXL $T=1564000 1214830 1 0 $X=1563998 $Y=1210890
X2145 15926 16463 16403 15687 15692 14586 16372 25 26 16293 SDFFNSRXL $T=1575960 1170550 0 180 $X=1564000 $Y=1166610
X2146 15937 16509 16504 15687 584 14691 16287 25 26 16417 SDFFNSRXL $T=1575960 1207450 0 180 $X=1564000 $Y=1203510
X2147 15942 16387 16484 16011 584 14466 16320 25 26 16418 SDFFNSRXL $T=1575960 1273870 0 180 $X=1564000 $Y=1269930
X2148 15941 16496 16503 595 15996 14671 16347 25 26 16394 SDFFNSRXL $T=1575960 1303390 1 180 $X=1564000 $Y=1303138
X2149 15926 16390 16508 15687 584 14623 16429 25 26 16368 SDFFNSRXL $T=1576420 1185310 1 180 $X=1564460 $Y=1185058
X2150 15942 16418 16481 16011 15692 14581 16441 25 26 16393 SDFFNSRXL $T=1569980 1273870 0 0 $X=1569978 $Y=1273618
X2151 8834 26 8814 8745 25 NOR2X1 $T=1059840 1104130 1 180 $X=1058460 $Y=1103878
X2152 8835 26 8860 8884 25 NOR2X1 $T=1058920 1177930 1 0 $X=1058918 $Y=1173990
X2153 8745 26 8945 8923 25 NOR2X1 $T=1064900 1104130 1 0 $X=1064898 $Y=1100190
X2154 8964 26 8816 8945 25 NOR2X1 $T=1069040 1111510 1 0 $X=1069038 $Y=1107570
X2155 9008 26 9014 9048 25 NOR2X1 $T=1070420 1081990 0 0 $X=1070418 $Y=1081738
X2156 9100 26 9079 9042 25 NOR2X1 $T=1076860 1089370 0 180 $X=1075480 $Y=1085430
X2157 9061 26 8749 9085 25 NOR2X1 $T=1076400 1104130 1 0 $X=1076398 $Y=1100190
X2158 9153 26 9085 9127 25 NOR2X1 $T=1077780 1096750 1 180 $X=1076400 $Y=1096498
X2159 8917 26 8742 9008 25 NOR2X1 $T=1081920 1074610 1 0 $X=1081918 $Y=1070670
X2160 9232 26 9219 9116 25 NOR2X1 $T=1085140 1089370 0 180 $X=1083760 $Y=1085430
X2161 9138 26 8961 9153 25 NOR2X1 $T=1087900 1104130 1 0 $X=1087898 $Y=1100190
X2162 8793 26 9282 9271 25 NOR2X1 $T=1088360 1148410 1 0 $X=1088358 $Y=1144470
X2163 8834 26 8870 9249 25 NOR2X1 $T=1092960 1074610 0 0 $X=1092958 $Y=1074358
X2164 9249 26 9352 9324 25 NOR2X1 $T=1093420 1067230 1 0 $X=1093418 $Y=1063290
X2165 9258 26 9101 9355 25 NOR2X1 $T=1093880 1089370 0 0 $X=1093878 $Y=1089118
X2166 9355 26 9362 9203 25 NOR2X1 $T=1095260 1096750 1 180 $X=1093880 $Y=1096498
X2167 9401 26 9327 9520 25 NOR2X1 $T=1096180 1045090 1 180 $X=1094800 $Y=1044838
X2168 8917 26 8822 9401 25 NOR2X1 $T=1095260 1059850 1 0 $X=1095258 $Y=1055910
X2169 8792 26 9415 9432 25 NOR2X1 $T=1097100 1148410 1 0 $X=1097098 $Y=1144470
X2170 8964 26 8931 9352 25 NOR2X1 $T=1097560 1074610 0 0 $X=1097558 $Y=1074358
X2171 9512 26 9228 9475 25 NOR2X1 $T=1098940 1074610 0 180 $X=1097560 $Y=1070670
X2172 9505 26 9475 9427 25 NOR2X1 $T=1101240 1081990 0 0 $X=1101238 $Y=1081738
X2173 9238 26 9003 9362 25 NOR2X1 $T=1101240 1104130 0 0 $X=1101238 $Y=1103878
X2174 9534 26 9102 9505 25 NOR2X1 $T=1105840 1081990 0 0 $X=1105838 $Y=1081738
X2175 9061 26 8880 9596 25 NOR2X1 $T=1109520 1074610 1 0 $X=1109518 $Y=1070670
X2176 9138 26 9005 9688 25 NOR2X1 $T=1109980 1074610 0 0 $X=1109978 $Y=1074358
X2177 9688 26 9596 9726 25 NOR2X1 $T=1110440 1067230 1 0 $X=1110438 $Y=1063290
X2178 9777 26 9196 9544 25 NOR2X1 $T=1111820 1096750 1 180 $X=1110440 $Y=1096498
X2179 9258 26 9243 9752 25 NOR2X1 $T=1110900 1059850 0 0 $X=1110898 $Y=1059598
X2180 9238 26 8980 9784 25 NOR2X1 $T=1114120 1074610 0 0 $X=1114118 $Y=1074358
X2181 9752 26 9784 9772 25 NOR2X1 $T=1114580 1059850 1 0 $X=1114578 $Y=1055910
X2182 9858 26 9785 9477 25 NOR2X1 $T=1115960 1081990 0 180 $X=1114580 $Y=1078050
X2183 9893 26 9715 9829 25 NOR2X1 $T=1118720 1045090 0 180 $X=1117340 $Y=1041150
X2184 9806 26 9270 9785 25 NOR2X1 $T=1119180 1081990 1 0 $X=1119178 $Y=1078050
X2185 10017 26 9916 9805 25 NOR2X1 $T=1122860 1096750 1 180 $X=1121480 $Y=1096498
X2186 10037 26 9916 9598 25 NOR2X1 $T=1122860 1104130 0 180 $X=1121480 $Y=1100190
X2187 10154 26 9916 9728 25 NOR2X1 $T=1129300 1104130 0 180 $X=1127920 $Y=1100190
X2188 10120 26 9196 9665 25 NOR2X1 $T=1129300 1170550 1 180 $X=1127920 $Y=1170298
X2189 10173 26 9916 9774 25 NOR2X1 $T=1129760 1104130 1 180 $X=1128380 $Y=1103878
X2190 10181 26 9916 9543 25 NOR2X1 $T=1130680 1118890 0 180 $X=1129300 $Y=1114950
X2191 10190 26 9916 10024 25 NOR2X1 $T=1132520 1096750 1 180 $X=1131140 $Y=1096498
X2192 10208 26 9916 9542 25 NOR2X1 $T=1132980 1111510 1 180 $X=1131600 $Y=1111258
X2193 10319 26 9916 9376 25 NOR2X1 $T=1138500 1126270 0 180 $X=1137120 $Y=1122330
X2194 10400 26 9196 9625 25 NOR2X1 $T=1140340 1163170 0 180 $X=1138960 $Y=1159230
X2195 10336 26 10294 10201 25 NOR2X1 $T=1140800 1045090 0 180 $X=1139420 $Y=1041150
X2196 9534 26 9518 10336 25 NOR2X1 $T=1139880 1059850 1 0 $X=1139878 $Y=1055910
X2197 9512 26 9437 10294 25 NOR2X1 $T=1139880 1059850 0 0 $X=1139878 $Y=1059598
X2198 10388 26 9916 10056 25 NOR2X1 $T=1141260 1111510 0 180 $X=1139880 $Y=1107570
X2199 10371 26 9916 10324 25 NOR2X1 $T=1142180 1126270 0 180 $X=1140800 $Y=1122330
X2200 9652 26 115 10613 25 NOR2X1 $T=1150920 1347670 1 0 $X=1150918 $Y=1343730
X2201 10616 26 10595 9090 25 NOR2X1 $T=1155060 1177930 1 180 $X=1153680 $Y=1177678
X2202 10598 26 10573 10228 25 NOR2X1 $T=1154600 1045090 1 0 $X=1154598 $Y=1041150
X2203 9806 26 10602 10573 25 NOR2X1 $T=1154600 1052470 0 0 $X=1154598 $Y=1052218
X2204 10619 26 10605 9272 25 NOR2X1 $T=1156440 1163170 1 180 $X=1155060 $Y=1162918
X2205 10605 26 10595 9054 25 NOR2X1 $T=1155520 1170550 0 0 $X=1155518 $Y=1170298
X2206 10644 26 9916 10267 25 NOR2X1 $T=1156900 1118890 0 180 $X=1155520 $Y=1114950
X2207 10619 26 10616 9049 25 NOR2X1 $T=1156900 1170550 0 180 $X=1155520 $Y=1166610
X2208 10646 26 9196 10630 25 NOR2X1 $T=1158280 1126270 1 180 $X=1156900 $Y=1126018
X2209 10717 26 134 10879 25 NOR2X1 $T=1162880 1318150 0 0 $X=1162878 $Y=1317898
X2210 10760 26 134 10906 25 NOR2X1 $T=1166560 1325530 1 0 $X=1166558 $Y=1321590
X2211 142 26 10880 10920 25 NOR2X1 $T=1169780 1347670 0 180 $X=1168400 $Y=1343730
X2212 10759 26 134 144 25 NOR2X1 $T=1168860 1347670 0 0 $X=1168858 $Y=1347418
X2213 10884 26 134 10934 25 NOR2X1 $T=1170700 1325530 1 0 $X=1170698 $Y=1321590
X2214 10983 26 10920 11081 25 NOR2X1 $T=1175300 1347670 0 180 $X=1173920 $Y=1343730
X2215 10975 26 134 11072 25 NOR2X1 $T=1174840 1325530 1 0 $X=1174838 $Y=1321590
X2216 153 26 10982 10983 25 NOR2X1 $T=1174840 1340290 1 0 $X=1174838 $Y=1336350
X2217 151 26 10934 11124 25 NOR2X1 $T=1178980 1325530 0 0 $X=1178978 $Y=1325278
X2218 161 26 11072 11149 25 NOR2X1 $T=1180820 1325530 0 180 $X=1179440 $Y=1321590
X2219 11011 26 11132 11150 25 NOR2X1 $T=1181280 1340290 0 0 $X=1181278 $Y=1340038
X2220 11124 26 11149 11189 25 NOR2X1 $T=1182200 1332910 1 0 $X=1182198 $Y=1328970
X2221 11124 26 11166 11164 25 NOR2X1 $T=1183120 1325530 0 0 $X=1183118 $Y=1325278
X2222 11422 26 11411 11391 25 NOR2X1 $T=1197840 1325530 1 180 $X=1196460 $Y=1325278
X2223 11428 26 9196 11498 25 NOR2X1 $T=1198300 1081990 1 180 $X=1196920 $Y=1081738
X2224 182 26 10879 11411 25 NOR2X1 $T=1199220 1318150 0 0 $X=1199218 $Y=1317898
X2225 11456 26 11254 11564 25 NOR2X1 $T=1201980 1340290 0 0 $X=1201978 $Y=1340038
X2226 187 26 10906 11422 25 NOR2X1 $T=1203820 1318150 1 180 $X=1202440 $Y=1317898
X2227 11749 26 11732 11848 25 NOR2X1 $T=1218540 1111510 0 180 $X=1217160 $Y=1107570
X2228 11786 26 207 11741 25 NOR2X1 $T=1218540 1347670 1 0 $X=1218538 $Y=1343730
X2229 11546 26 11561 11862 25 NOR2X1 $T=1219460 1185310 0 0 $X=1219458 $Y=1185058
X2230 211 26 11899 207 25 NOR2X1 $T=1221760 1340290 0 180 $X=1220380 $Y=1336350
X2231 11926 26 11147 11749 25 NOR2X1 $T=1221300 1111510 0 0 $X=1221298 $Y=1111258
X2232 11941 26 11437 11732 25 NOR2X1 $T=1222680 1111510 0 180 $X=1221300 $Y=1107570
X2233 11901 26 10967 11798 25 NOR2X1 $T=1222680 1126270 0 0 $X=1222678 $Y=1126018
X2234 212 26 10876 11786 25 NOR2X1 $T=1224060 1347670 0 180 $X=1222680 $Y=1343730
X2235 11901 26 11449 11984 25 NOR2X1 $T=1224520 1170550 0 0 $X=1224518 $Y=1170298
X2236 12190 26 12078 221 25 NOR2X1 $T=1230500 1296010 1 180 $X=1229120 $Y=1295758
X2237 11941 26 11425 12219 25 NOR2X1 $T=1233720 1170550 0 0 $X=1233718 $Y=1170298
X2238 11926 26 11314 12249 25 NOR2X1 $T=1234640 1163170 1 0 $X=1234638 $Y=1159230
X2239 12253 26 11322 12223 25 NOR2X1 $T=1237860 1104130 0 0 $X=1237858 $Y=1103878
X2240 12278 26 12266 12152 25 NOR2X1 $T=1239700 1111510 0 180 $X=1238320 $Y=1107570
X2241 12333 26 12223 12161 25 NOR2X1 $T=1240620 1104130 0 180 $X=1239240 $Y=1100190
X2242 12249 26 12219 12347 25 NOR2X1 $T=1241540 1170550 1 0 $X=1241538 $Y=1166610
X2243 11112 26 11242 12390 25 NOR2X1 $T=1243840 1052470 1 0 $X=1243838 $Y=1048530
X2244 11363 26 11242 12451 25 NOR2X1 $T=1243840 1081990 0 0 $X=1243838 $Y=1081738
X2245 12393 26 11323 12266 25 NOR2X1 $T=1248900 1118890 0 0 $X=1248898 $Y=1118638
X2246 12551 26 12539 12512 25 NOR2X1 $T=1251660 1081990 1 180 $X=1250280 $Y=1081738
X2247 12582 26 11063 12464 25 NOR2X1 $T=1252120 1059850 1 0 $X=1252118 $Y=1055910
X2248 12500 26 11275 12333 25 NOR2X1 $T=1253500 1104130 0 0 $X=1253498 $Y=1103878
X2249 12704 26 12464 12594 25 NOR2X1 $T=1258100 1059850 0 180 $X=1256720 $Y=1055910
X2250 12762 26 12706 12453 25 NOR2X1 $T=1259480 1067230 1 180 $X=1258100 $Y=1066978
X2251 12685 26 11066 12704 25 NOR2X1 $T=1260860 1059850 0 0 $X=1260858 $Y=1059598
X2252 12814 26 11344 12691 25 NOR2X1 $T=1262240 1096750 0 180 $X=1260860 $Y=1092810
X2253 12857 26 11087 12762 25 NOR2X1 $T=1271440 1074610 1 0 $X=1271438 $Y=1070670
X2254 12943 26 11243 12880 25 NOR2X1 $T=1273280 1089370 1 180 $X=1271900 $Y=1089118
X2255 12929 26 11421 13058 25 NOR2X1 $T=1273280 1111510 1 0 $X=1273278 $Y=1107570
X2256 13058 26 13030 12988 25 NOR2X1 $T=1274660 1104130 1 0 $X=1274658 $Y=1100190
X2257 12685 26 12889 13054 25 NOR2X1 $T=1277880 1067230 1 0 $X=1277878 $Y=1063290
X2258 13252 26 13248 13165 25 NOR2X1 $T=1284320 1170550 0 180 $X=1282940 $Y=1166610
X2259 12814 26 12874 13372 25 NOR2X1 $T=1283860 1096750 1 0 $X=1283858 $Y=1092810
X2260 12857 26 12744 13251 25 NOR2X1 $T=1284780 1081990 1 0 $X=1284778 $Y=1078050
X2261 13054 26 13297 13381 25 NOR2X1 $T=1285240 1059850 0 0 $X=1285238 $Y=1059598
X2262 13251 26 13307 13324 25 NOR2X1 $T=1285700 1074610 1 0 $X=1285698 $Y=1070670
X2263 12834 26 12729 13362 25 NOR2X1 $T=1286160 1104130 0 0 $X=1286158 $Y=1103878
X2264 12730 26 12926 13307 25 NOR2X1 $T=1288920 1081990 0 0 $X=1288918 $Y=1081738
X2265 12943 26 12927 13389 25 NOR2X1 $T=1288920 1096750 0 0 $X=1288918 $Y=1096498
X2266 12582 26 13161 13297 25 NOR2X1 $T=1289840 1059850 1 0 $X=1289838 $Y=1055910
X2267 13389 26 13372 13393 25 NOR2X1 $T=1289840 1089370 0 0 $X=1289838 $Y=1089118
X2268 12500 26 12463 13448 25 NOR2X1 $T=1292140 1126270 1 0 $X=1292138 $Y=1122330
X2269 13440 26 13446 13451 25 NOR2X1 $T=1292600 1067230 0 0 $X=1292598 $Y=1066978
X2270 12393 26 11177 13501 25 NOR2X1 $T=1293060 1141030 0 0 $X=1293058 $Y=1140778
X2271 12929 26 13453 13506 25 NOR2X1 $T=1295820 1111510 1 0 $X=1295818 $Y=1107570
X2272 12253 26 11345 13582 25 NOR2X1 $T=1296740 1126270 1 0 $X=1296738 $Y=1122330
X2273 13506 26 13362 13546 25 NOR2X1 $T=1297200 1104130 0 0 $X=1297198 $Y=1103878
X2274 13448 26 13582 13631 25 NOR2X1 $T=1300420 1126270 1 0 $X=1300418 $Y=1122330
X2275 13554 26 13501 13651 25 NOR2X1 $T=1303180 1141030 1 0 $X=1303178 $Y=1137090
X2276 15933 26 368 15952 25 NOR2X1 $T=1526740 1170550 1 180 $X=1525360 $Y=1170298
X2277 558 26 15949 15939 25 NOR2X1 $T=1526740 1200070 0 180 $X=1525360 $Y=1196130
X2278 15986 26 15952 15944 25 NOR2X1 $T=1527200 1177930 0 180 $X=1525820 $Y=1173990
X2279 13915 26 375 15980 25 NOR2X1 $T=1527200 1259110 0 0 $X=1527198 $Y=1258858
X2280 15977 26 416 16051 25 NOR2X1 $T=1528580 1192690 0 180 $X=1527200 $Y=1188750
X2281 561 26 378 15986 25 NOR2X1 $T=1530880 1177930 1 180 $X=1529500 $Y=1177678
X2282 15933 26 369 16040 25 NOR2X1 $T=1531800 1177930 1 0 $X=1531798 $Y=1173990
X2283 16032 26 16028 16026 25 NOR2X1 $T=1533180 1332910 1 180 $X=1531800 $Y=1332658
X2284 415 26 16035 16042 25 NOR2X1 $T=1532720 1303390 0 0 $X=1532718 $Y=1303138
X2285 16073 26 16033 15955 25 NOR2X1 $T=1534100 1155790 1 180 $X=1532720 $Y=1155538
X2286 521 26 389 16050 25 NOR2X1 $T=1533180 1185310 1 0 $X=1533178 $Y=1181370
X2287 16047 26 16040 16085 25 NOR2X1 $T=1535020 1177930 1 180 $X=1533640 $Y=1177678
X2288 564 26 373 16047 25 NOR2X1 $T=1535940 1251730 0 180 $X=1534560 $Y=1247790
X2289 15980 26 16059 15973 25 NOR2X1 $T=1535940 1251730 0 0 $X=1535938 $Y=1251478
X2290 521 26 386 16060 25 NOR2X1 $T=1535940 1259110 0 0 $X=1535938 $Y=1258858
X2291 16070 26 16051 16056 25 NOR2X1 $T=1537320 1192690 0 180 $X=1535940 $Y=1188750
X2292 566 26 16061 15781 25 NOR2X1 $T=1537320 1296010 0 180 $X=1535940 $Y=1292070
X2293 16050 26 16066 16067 25 NOR2X1 $T=1536400 1163170 0 0 $X=1536398 $Y=1162918
X2294 558 26 16065 16127 25 NOR2X1 $T=1536400 1207450 0 0 $X=1536398 $Y=1207198
X2295 561 26 398 16077 25 NOR2X1 $T=1536400 1236970 1 0 $X=1536398 $Y=1233030
X2296 16047 26 16068 16123 25 NOR2X1 $T=1536400 1244350 1 0 $X=1536398 $Y=1240410
X2297 16042 26 16050 15945 25 NOR2X1 $T=1536400 1303390 1 0 $X=1536398 $Y=1299450
X2298 16074 26 386 16065 25 NOR2X1 $T=1537780 1207450 0 180 $X=1536400 $Y=1203510
X2299 16100 26 550 16028 25 NOR2X1 $T=1537780 1340290 0 180 $X=1536400 $Y=1336350
X2300 561 26 375 16078 25 NOR2X1 $T=1537320 1177930 1 0 $X=1537318 $Y=1173990
X2301 567 26 364 16086 25 NOR2X1 $T=1538700 1273870 1 180 $X=1537320 $Y=1273618
X2302 16095 26 535 16032 25 NOR2X1 $T=1538700 1332910 1 180 $X=1537320 $Y=1332658
X2303 15981 26 415 16066 25 NOR2X1 $T=1537780 1148410 1 0 $X=1537778 $Y=1144470
X2304 521 26 369 16073 25 NOR2X1 $T=1537780 1155790 0 0 $X=1537778 $Y=1155538
X2305 16078 26 16087 16158 25 NOR2X1 $T=1537780 1170550 0 0 $X=1537778 $Y=1170298
X2306 16060 26 16093 16034 25 NOR2X1 $T=1537780 1259110 1 0 $X=1537778 $Y=1255170
X2307 16035 26 458 16118 25 NOR2X1 $T=1537780 1303390 0 0 $X=1537778 $Y=1303138
X2308 15983 26 388 16151 25 NOR2X1 $T=1538240 1214830 0 0 $X=1538238 $Y=1214578
X2309 375 26 16099 16059 25 NOR2X1 $T=1538240 1251730 1 0 $X=1538238 $Y=1247790
X2310 16072 26 412 16033 25 NOR2X1 $T=1538700 1148410 0 0 $X=1538698 $Y=1148158
X2311 16072 26 398 16087 25 NOR2X1 $T=1538700 1163170 1 0 $X=1538698 $Y=1159230
X2312 16086 26 16104 16069 25 NOR2X1 $T=1538700 1273870 1 0 $X=1538698 $Y=1269930
X2313 16100 26 485 16154 25 NOR2X1 $T=1538700 1340290 1 0 $X=1538698 $Y=1336350
X2314 16099 26 13974 16093 25 NOR2X1 $T=1540080 1259110 1 0 $X=1540078 $Y=1255170
X2315 15934 26 370 16162 25 NOR2X1 $T=1541000 1318150 0 0 $X=1540998 $Y=1317898
X2316 16130 26 373 16061 25 NOR2X1 $T=1542380 1296010 0 180 $X=1541000 $Y=1292070
X2317 16077 26 16157 16152 25 NOR2X1 $T=1541920 1236970 1 0 $X=1541918 $Y=1233030
X2318 16163 26 16155 16169 25 NOR2X1 $T=1543300 1155790 1 180 $X=1541920 $Y=1155538
X2319 574 26 16151 16192 25 NOR2X1 $T=1543300 1222210 0 180 $X=1541920 $Y=1218270
X2320 16078 26 16166 16216 25 NOR2X1 $T=1542380 1214830 1 0 $X=1542378 $Y=1210890
X2321 571 26 16167 16195 25 NOR2X1 $T=1542380 1251730 1 0 $X=1542378 $Y=1247790
X2322 570 26 16162 16094 25 NOR2X1 $T=1542380 1325530 1 0 $X=1542378 $Y=1321590
X2323 570 26 16154 16126 25 NOR2X1 $T=1542380 1340290 1 0 $X=1542378 $Y=1336350
X2324 16163 26 16165 16156 25 NOR2X1 $T=1543760 1200070 1 180 $X=1542380 $Y=1199818
X2325 16208 26 375 16104 25 NOR2X1 $T=1543760 1273870 0 180 $X=1542380 $Y=1269930
X2326 15983 26 458 16166 25 NOR2X1 $T=1542840 1214830 0 0 $X=1542838 $Y=1214578
X2327 15934 26 535 16179 25 NOR2X1 $T=1542840 1318150 0 0 $X=1542838 $Y=1317898
X2328 575 26 16118 16225 25 NOR2X1 $T=1544220 1303390 1 180 $X=1542840 $Y=1303138
X2329 561 26 370 16070 25 NOR2X1 $T=1543300 1192690 1 0 $X=1543298 $Y=1188750
X2330 521 26 415 16219 25 NOR2X1 $T=1543300 1266490 0 0 $X=1543298 $Y=1266238
X2331 561 26 364 16163 25 NOR2X1 $T=1543760 1170550 1 0 $X=1543758 $Y=1166610
X2332 364 26 16130 16196 25 NOR2X1 $T=1543760 1288630 0 0 $X=1543758 $Y=1288378
X2333 16074 26 401 16165 25 NOR2X1 $T=1544220 1207450 1 0 $X=1544218 $Y=1203510
X2334 16201 26 388 16068 25 NOR2X1 $T=1545600 1244350 1 180 $X=1544220 $Y=1244098
X2335 16187 26 389 16286 25 NOR2X1 $T=1544680 1155790 1 0 $X=1544678 $Y=1151850
X2336 575 26 16196 16181 25 NOR2X1 $T=1546060 1296010 0 180 $X=1544680 $Y=1292070
X2337 16177 26 398 16157 25 NOR2X1 $T=1545140 1236970 1 0 $X=1545138 $Y=1233030
X2338 16187 26 378 16229 25 NOR2X1 $T=1545600 1155790 0 0 $X=1545598 $Y=1155538
X2339 16201 26 378 16167 25 NOR2X1 $T=1546060 1251730 1 0 $X=1546058 $Y=1247790
X2340 16208 26 386 16255 25 NOR2X1 $T=1546060 1273870 1 0 $X=1546058 $Y=1269930
X2341 583 26 16179 15893 25 NOR2X1 $T=1547440 1325530 0 180 $X=1546060 $Y=1321590
X2342 16177 26 13974 16269 25 NOR2X1 $T=1548360 1236970 1 0 $X=1548358 $Y=1233030
X2343 521 26 13974 16268 25 NOR2X1 $T=1549280 1155790 0 0 $X=1549278 $Y=1155538
X2344 585 26 16255 16251 25 NOR2X1 $T=1550200 1273870 1 0 $X=1550198 $Y=1269930
X2345 16219 26 16271 16296 25 NOR2X1 $T=1550200 1281250 1 0 $X=1550198 $Y=1277310
X2346 585 26 16269 16275 25 NOR2X1 $T=1550660 1236970 0 0 $X=1550658 $Y=1236718
X2347 561 26 485 16292 25 NOR2X1 $T=1552500 1155790 0 0 $X=1552498 $Y=1155538
X2348 588 26 16291 16270 25 NOR2X1 $T=1552960 1170550 0 0 $X=1552958 $Y=1170298
X2349 16268 26 16286 16338 25 NOR2X1 $T=1553420 1155790 1 0 $X=1553418 $Y=1151850
X2350 16219 26 16306 16314 25 NOR2X1 $T=1554800 1192690 1 0 $X=1554798 $Y=1188750
X2351 16313 26 389 16306 25 NOR2X1 $T=1556180 1170550 0 180 $X=1554800 $Y=1166610
X2352 16363 26 389 16271 25 NOR2X1 $T=1556640 1281250 0 180 $X=1555260 $Y=1277310
X2353 16292 26 16229 16365 25 NOR2X1 $T=1556180 1155790 0 0 $X=1556178 $Y=1155538
X2354 16313 26 485 16291 25 NOR2X1 $T=1556180 1170550 0 0 $X=1556178 $Y=1170298
X2355 16363 26 368 16373 25 NOR2X1 $T=1560320 1281250 1 180 $X=1558940 $Y=1280998
X2356 561 26 416 588 25 NOR2X1 $T=1559860 1177930 1 0 $X=1559858 $Y=1173990
X2357 593 26 16373 16327 25 NOR2X1 $T=1560320 1288630 1 0 $X=1560318 $Y=1284690
X2358 8677 25 26 8734 CLKINVX1 $T=1040060 1155790 1 0 $X=1040058 $Y=1151850
X2359 8734 25 26 8738 CLKINVX1 $T=1043740 1148410 1 0 $X=1043738 $Y=1144470
X2360 8737 25 26 8818 CLKINVX1 $T=1044660 1141030 0 180 $X=1043740 $Y=1137090
X2361 8742 25 26 8822 CLKINVX1 $T=1045120 1133650 1 180 $X=1044200 $Y=1133398
X2362 8741 25 26 8737 CLKINVX1 $T=1045120 1141030 1 180 $X=1044200 $Y=1140778
X2363 8745 25 26 8882 CLKINVX1 $T=1047420 1111510 0 180 $X=1046500 $Y=1107570
X2364 8750 25 26 8819 CLKINVX1 $T=1052480 1148410 1 0 $X=1052478 $Y=1144470
X2365 8749 25 26 8880 CLKINVX1 $T=1058460 1148410 1 0 $X=1058458 $Y=1144470
X2366 8859 25 26 8750 CLKINVX1 $T=1059840 1148410 1 180 $X=1058920 $Y=1148158
X2367 8920 25 26 8743 CLKINVX1 $T=1059840 1155790 1 180 $X=1058920 $Y=1155538
X2368 8932 25 26 8835 CLKINVX1 $T=1059840 1177930 1 180 $X=1058920 $Y=1177678
X2369 8858 25 26 8877 CLKINVX1 $T=1059380 1081990 0 0 $X=1059378 $Y=1081738
X2370 8736 25 26 8881 CLKINVX1 $T=1059380 1192690 0 0 $X=1059378 $Y=1192438
X2371 8946 25 26 8838 CLKINVX1 $T=1061220 1163170 1 180 $X=1060300 $Y=1162918
X2372 8872 25 26 8733 CLKINVX1 $T=1061220 1170550 1 180 $X=1060300 $Y=1170298
X2373 8943 25 26 8793 CLKINVX1 $T=1063060 1148410 0 180 $X=1062140 $Y=1144470
X2374 8883 25 26 8948 CLKINVX1 $T=1064440 1192690 0 0 $X=1064438 $Y=1192438
X2375 8860 25 26 8954 CLKINVX1 $T=1064900 1185310 1 0 $X=1064898 $Y=1181370
X2376 8792 25 26 8975 CLKINVX1 $T=1066280 1148410 1 0 $X=1066278 $Y=1144470
X2377 9042 25 26 8913 CLKINVX1 $T=1070880 1096750 0 180 $X=1069960 $Y=1092810
X2378 9075 25 26 9137 CLKINVX1 $T=1075480 1192690 0 0 $X=1075478 $Y=1192438
X2379 8824 25 26 8976 CLKINVX1 $T=1076400 1133650 1 0 $X=1076398 $Y=1129710
X2380 9081 25 26 9129 CLKINVX1 $T=1077320 1200070 1 0 $X=1077318 $Y=1196130
X2381 9110 25 26 9114 CLKINVX1 $T=1077780 1059850 0 0 $X=1077778 $Y=1059598
X2382 9119 25 26 8935 CLKINVX1 $T=1077780 1148410 0 0 $X=1077778 $Y=1148158
X2383 9177 25 26 8824 CLKINVX1 $T=1078700 1133650 1 180 $X=1077780 $Y=1133398
X2384 9253 25 26 9094 CLKINVX1 $T=1083760 1222210 0 180 $X=1082840 $Y=1218270
X2385 9141 25 26 8792 CLKINVX1 $T=1083300 1148410 1 0 $X=1083298 $Y=1144470
X2386 9232 25 26 9254 CLKINVX1 $T=1086980 1081990 0 0 $X=1086978 $Y=1081738
X2387 8732 25 26 9225 CLKINVX1 $T=1086980 1185310 0 0 $X=1086978 $Y=1185058
X2388 9220 25 26 9290 CLKINVX1 $T=1088820 1089370 0 0 $X=1088818 $Y=1089118
X2389 9327 25 26 9338 CLKINVX1 $T=1092500 1052470 0 0 $X=1092498 $Y=1052218
X2390 9325 25 26 9377 CLKINVX1 $T=1092500 1185310 0 0 $X=1092498 $Y=1185058
X2391 9250 25 26 9199 CLKINVX1 $T=1092960 1081990 0 0 $X=1092958 $Y=1081738
X2392 9328 25 26 9420 CLKINVX1 $T=1092960 1229590 0 0 $X=1092958 $Y=1229338
X2393 9395 25 26 9329 CLKINVX1 $T=1093880 1266490 1 180 $X=1092960 $Y=1266238
X2394 9340 25 26 9316 CLKINVX1 $T=1093880 1273870 0 180 $X=1092960 $Y=1269930
X2395 9128 25 26 9393 CLKINVX1 $T=1093420 1177930 1 0 $X=1093418 $Y=1173990
X2396 9353 25 26 9013 CLKINVX1 $T=1093880 1170550 0 0 $X=1093878 $Y=1170298
X2397 9300 25 26 9403 CLKINVX1 $T=1093880 1192690 0 0 $X=1093878 $Y=1192438
X2398 9335 25 26 9343 CLKINVX1 $T=1094800 1214830 1 180 $X=1093880 $Y=1214578
X2399 9359 25 26 8952 CLKINVX1 $T=1096180 1133650 1 180 $X=1095260 $Y=1133398
X2400 9419 25 26 48 CLKINVX1 $T=1096180 1340290 1 180 $X=1095260 $Y=1340038
X2401 9417 25 26 9350 CLKINVX1 $T=1097560 1251730 0 180 $X=1096640 $Y=1247790
X2402 9407 25 26 9344 CLKINVX1 $T=1097100 1229590 0 0 $X=1097098 $Y=1229338
X2403 9299 25 26 9281 CLKINVX1 $T=1099860 1089370 0 0 $X=1099858 $Y=1089118
X2404 9358 25 26 9379 CLKINVX1 $T=1099860 1163170 1 0 $X=1099858 $Y=1159230
X2405 9394 25 26 9354 CLKINVX1 $T=1099860 1222210 1 0 $X=1099858 $Y=1218270
X2406 9351 25 26 9488 CLKINVX1 $T=1099860 1251730 1 0 $X=1099858 $Y=1247790
X2407 9505 25 26 9563 CLKINVX1 $T=1100780 1089370 0 180 $X=1099860 $Y=1085430
X2408 9547 25 26 9668 CLKINVX1 $T=1103540 1303390 1 0 $X=1103538 $Y=1299450
X2409 9471 25 26 9248 CLKINVX1 $T=1104920 1059850 0 180 $X=1104000 $Y=1055910
X2410 9559 25 26 9438 CLKINVX1 $T=1104460 1244350 1 0 $X=1104458 $Y=1240410
X2411 9541 25 26 9549 CLKINVX1 $T=1104920 1207450 0 0 $X=1104918 $Y=1207198
X2412 9576 25 26 9426 CLKINVX1 $T=1104920 1288630 0 0 $X=1104918 $Y=1288378
X2413 9425 25 26 9651 CLKINVX1 $T=1106300 1259110 0 0 $X=1106298 $Y=1258858
X2414 9681 25 26 9436 CLKINVX1 $T=1111360 1244350 1 180 $X=1110440 $Y=1244098
X2415 9487 25 26 9791 CLKINVX1 $T=1110900 1170550 0 0 $X=1110898 $Y=1170298
X2416 9903 25 26 46 CLKINVX1 $T=1111820 1288630 1 180 $X=1110900 $Y=1288378
X2417 72 25 26 9687 CLKINVX1 $T=1111820 1310770 0 180 $X=1110900 $Y=1306830
X2418 9748 25 26 9531 CLKINVX1 $T=1113660 1200070 1 180 $X=1112740 $Y=1199818
X2419 9594 25 26 9803 CLKINVX1 $T=1113660 1296010 1 0 $X=1113658 $Y=1292070
X2420 9753 25 26 9807 CLKINVX1 $T=1115500 1200070 0 0 $X=1115498 $Y=1199818
X2421 9744 25 26 9827 CLKINVX1 $T=1115500 1266490 1 0 $X=1115498 $Y=1262550
X2422 9814 25 26 9800 CLKINVX1 $T=1116420 1236970 1 0 $X=1116418 $Y=1233030
X2423 9382 25 26 44 CLKINVX1 $T=1116880 1214830 1 0 $X=1116878 $Y=1210890
X2424 77 25 26 9871 CLKINVX1 $T=1116880 1318150 0 0 $X=1116878 $Y=1317898
X2425 9768 25 26 9746 CLKINVX1 $T=1117800 1281250 0 0 $X=1117798 $Y=1280998
X2426 9667 25 26 9570 CLKINVX1 $T=1120560 1163170 1 0 $X=1120558 $Y=1159230
X2427 9849 25 26 9862 CLKINVX1 $T=1122860 1045090 0 0 $X=1122858 $Y=1044838
X2428 9978 25 26 9927 CLKINVX1 $T=1124700 1081990 0 180 $X=1123780 $Y=1078050
X2429 9930 25 26 9915 CLKINVX1 $T=1127460 1310770 1 0 $X=1127458 $Y=1306830
X2430 10052 25 26 10051 CLKINVX1 $T=1128380 1288630 1 180 $X=1127460 $Y=1288378
X2431 98 25 26 10047 CLKINVX1 $T=1128380 1303390 0 180 $X=1127460 $Y=1299450
X2432 9858 25 26 9904 CLKINVX1 $T=1127920 1081990 1 0 $X=1127918 $Y=1078050
X2433 81 25 26 10166 CLKINVX1 $T=1130680 1303390 1 0 $X=1130678 $Y=1299450
X2434 10139 25 26 10110 CLKINVX1 $T=1132520 1288630 0 180 $X=1131600 $Y=1284690
X2435 10080 25 26 10217 CLKINVX1 $T=1134360 1185310 0 0 $X=1134358 $Y=1185058
X2436 9372 25 26 10220 CLKINVX1 $T=1134360 1303390 1 0 $X=1134358 $Y=1299450
X2437 104 25 26 10274 CLKINVX1 $T=1137580 1303390 1 0 $X=1137578 $Y=1299450
X2438 10256 25 26 10404 CLKINVX1 $T=1138500 1340290 0 0 $X=1138498 $Y=1340038
X2439 10106 25 26 10322 CLKINVX1 $T=1139880 1118890 0 0 $X=1139878 $Y=1118638
X2440 107 25 26 10337 CLKINVX1 $T=1140340 1325530 0 0 $X=1140338 $Y=1325278
X2441 10017 25 26 10397 CLKINVX1 $T=1140800 1096750 0 0 $X=1140798 $Y=1096498
X2442 10337 25 26 10353 CLKINVX1 $T=1140800 1303390 1 0 $X=1140798 $Y=1299450
X2443 10407 25 26 10389 CLKINVX1 $T=1144480 1111510 0 180 $X=1143560 $Y=1107570
X2444 10390 25 26 10443 CLKINVX1 $T=1144020 1229590 1 0 $X=1144018 $Y=1225650
X2445 10173 25 26 10423 CLKINVX1 $T=1144480 1111510 1 0 $X=1144478 $Y=1107570
X2446 112 25 26 9924 CLKINVX1 $T=1144480 1318150 1 0 $X=1144478 $Y=1314210
X2447 9967 25 26 10485 CLKINVX1 $T=1144940 1281250 1 0 $X=1144938 $Y=1277310
X2448 10439 25 26 10418 CLKINVX1 $T=1146320 1185310 1 180 $X=1145400 $Y=1185058
X2449 10447 25 26 10399 CLKINVX1 $T=1148620 1089370 0 180 $X=1147700 $Y=1085430
X2450 10096 25 26 9725 CLKINVX1 $T=1149540 1045090 0 0 $X=1149538 $Y=1044838
X2451 10249 25 26 116 CLKINVX1 $T=1150460 1340290 0 0 $X=1150458 $Y=1340038
X2452 10545 25 26 10538 CLKINVX1 $T=1151840 1118890 1 180 $X=1150920 $Y=1118638
X2453 10469 25 26 10106 CLKINVX1 $T=1152300 1126270 1 180 $X=1151380 $Y=1126018
X2454 10548 25 26 10526 CLKINVX1 $T=1152760 1104130 0 180 $X=1151840 $Y=1100190
X2455 10335 25 26 121 CLKINVX1 $T=1153680 1340290 0 0 $X=1153678 $Y=1340038
X2456 10612 25 26 9913 CLKINVX1 $T=1155060 1296010 1 180 $X=1154140 $Y=1295758
X2457 10440 25 26 10717 CLKINVX1 $T=1155520 1310770 1 0 $X=1155518 $Y=1306830
X2458 10037 25 26 10653 CLKINVX1 $T=1157360 1104130 1 0 $X=1157358 $Y=1100190
X2459 10573 25 26 10744 CLKINVX1 $T=1157820 1037710 0 0 $X=1157818 $Y=1037458
X2460 10849 25 26 10102 CLKINVX1 $T=1158740 1281250 0 180 $X=1157820 $Y=1277310
X2461 10598 25 26 10732 CLKINVX1 $T=1158280 1045090 1 0 $X=1158278 $Y=1041150
X2462 10769 25 26 9928 CLKINVX1 $T=1159200 1296010 1 180 $X=1158280 $Y=1295758
X2463 10674 25 26 10555 CLKINVX1 $T=1159200 1303390 0 180 $X=1158280 $Y=1299450
X2464 10190 25 26 10728 CLKINVX1 $T=1159200 1096750 0 0 $X=1159198 $Y=1096498
X2465 10730 25 26 10121 CLKINVX1 $T=1161960 1236970 1 180 $X=1161040 $Y=1236718
X2466 129 25 26 10657 CLKINVX1 $T=1162420 1340290 1 180 $X=1161500 $Y=1340038
X2467 10486 25 26 10470 CLKINVX1 $T=1161960 1177930 1 0 $X=1161958 $Y=1173990
X2468 9729 25 26 9525 CLKINVX1 $T=1161960 1177930 0 0 $X=1161958 $Y=1177678
X2469 10714 25 26 10799 CLKINVX1 $T=1161960 1214830 0 0 $X=1161958 $Y=1214578
X2470 10737 25 26 10747 CLKINVX1 $T=1161960 1340290 1 0 $X=1161958 $Y=1336350
X2471 10149 25 26 10759 CLKINVX1 $T=1161960 1347670 0 0 $X=1161958 $Y=1347418
X2472 10624 25 26 10709 CLKINVX1 $T=1162880 1118890 0 180 $X=1161960 $Y=1114950
X2473 10851 25 26 10684 CLKINVX1 $T=1163340 1089370 0 180 $X=1162420 $Y=1085430
X2474 10437 25 26 10760 CLKINVX1 $T=1162880 1325530 1 0 $X=1162878 $Y=1321590
X2475 10736 25 26 10761 CLKINVX1 $T=1162880 1332910 1 0 $X=1162878 $Y=1328970
X2476 10488 25 26 10770 CLKINVX1 $T=1162880 1347670 1 0 $X=1162878 $Y=1343730
X2477 10800 25 26 10053 CLKINVX1 $T=1164720 1229590 1 180 $X=1163800 $Y=1229338
X2478 10781 25 26 10436 CLKINVX1 $T=1164720 1244350 1 180 $X=1163800 $Y=1244098
X2479 10589 25 26 10889 CLKINVX1 $T=1164260 1325530 0 0 $X=1164258 $Y=1325278
X2480 10683 25 26 10857 CLKINVX1 $T=1166100 1266490 0 0 $X=1166098 $Y=1266238
X2481 10843 25 26 10279 CLKINVX1 $T=1167480 1266490 0 180 $X=1166560 $Y=1262550
X2482 126 25 26 10486 CLKINVX1 $T=1167020 1177930 0 0 $X=1167018 $Y=1177678
X2483 10445 25 26 10869 CLKINVX1 $T=1167480 1273870 0 0 $X=1167478 $Y=1273618
X2484 140 25 26 10616 CLKINVX1 $T=1169320 1185310 0 180 $X=1168400 $Y=1181370
X2485 10842 25 26 10884 CLKINVX1 $T=1168860 1318150 0 0 $X=1168858 $Y=1317898
X2486 10522 25 26 10885 CLKINVX1 $T=1168860 1332910 0 0 $X=1168858 $Y=1332658
X2487 74 25 26 10924 CLKINVX1 $T=1169320 1288630 0 0 $X=1169318 $Y=1288378
X2488 9966 25 26 10942 CLKINVX1 $T=1169780 1266490 1 0 $X=1169778 $Y=1262550
X2489 10878 25 26 10948 CLKINVX1 $T=1171160 1177930 0 0 $X=1171158 $Y=1177678
X2490 9781 25 26 10999 CLKINVX1 $T=1172540 1251730 1 0 $X=1172538 $Y=1247790
X2491 11043 25 26 10743 CLKINVX1 $T=1173920 1310770 0 180 $X=1173000 $Y=1306830
X2492 10973 25 26 10566 CLKINVX1 $T=1174380 1251730 1 180 $X=1173460 $Y=1251478
X2493 10801 25 26 10975 CLKINVX1 $T=1174380 1318150 0 0 $X=1174378 $Y=1317898
X2494 10980 25 26 10929 CLKINVX1 $T=1175760 1089370 0 180 $X=1174840 $Y=1085430
X2495 141 25 26 10530 CLKINVX1 $T=1175300 1177930 0 0 $X=1175298 $Y=1177678
X2496 11007 25 26 10922 CLKINVX1 $T=1176220 1111510 1 180 $X=1175300 $Y=1111258
X2497 10269 25 26 11071 CLKINVX1 $T=1175760 1251730 1 0 $X=1175758 $Y=1247790
X2498 10983 25 26 11075 CLKINVX1 $T=1175760 1347670 0 0 $X=1175758 $Y=1347418
X2499 11086 25 26 10840 CLKINVX1 $T=1179900 1310770 1 180 $X=1178980 $Y=1310518
X2500 11124 25 26 11073 CLKINVX1 $T=1179900 1332910 1 180 $X=1178980 $Y=1332658
X2501 11084 25 26 11090 CLKINVX1 $T=1179440 1185310 0 0 $X=1179438 $Y=1185058
X2502 10927 25 26 11056 CLKINVX1 $T=1180360 1037710 1 180 $X=1179440 $Y=1037458
X2503 10955 25 26 11109 CLKINVX1 $T=1179900 1266490 1 0 $X=1179898 $Y=1262550
X2504 159 25 26 10809 CLKINVX1 $T=1181740 1318150 0 180 $X=1180820 $Y=1314210
X2505 10644 25 26 11128 CLKINVX1 $T=1182200 1104130 0 0 $X=1182198 $Y=1103878
X2506 11064 25 26 11139 CLKINVX1 $T=1182200 1332910 0 0 $X=1182198 $Y=1332658
X2507 11038 25 26 11205 CLKINVX1 $T=1183580 1037710 0 0 $X=1183578 $Y=1037458
X2508 11196 25 26 11172 CLKINVX1 $T=1185420 1133650 0 180 $X=1184500 $Y=1129710
X2509 11197 25 26 11203 CLKINVX1 $T=1184960 1148410 1 0 $X=1184958 $Y=1144470
X2510 10945 25 26 11236 CLKINVX1 $T=1185880 1104130 1 0 $X=1185878 $Y=1100190
X2511 11143 25 26 11235 CLKINVX1 $T=1186340 1096750 1 0 $X=1186338 $Y=1092810
X2512 173 25 26 10595 CLKINVX1 $T=1187720 1185310 0 180 $X=1186800 $Y=1181370
X2513 10994 25 26 11153 CLKINVX1 $T=1188180 1059850 1 180 $X=1187260 $Y=1059598
X2514 11282 25 26 9965 CLKINVX1 $T=1188640 1259110 1 180 $X=1187720 $Y=1258858
X2515 11138 25 26 11351 CLKINVX1 $T=1192320 1059850 0 0 $X=1192318 $Y=1059598
X2516 11166 25 26 11334 CLKINVX1 $T=1192780 1325530 1 0 $X=1192778 $Y=1321590
X2517 11219 25 26 11308 CLKINVX1 $T=1194160 1118890 0 180 $X=1193240 $Y=1114950
X2518 11415 25 26 10289 CLKINVX1 $T=1196460 1200070 0 180 $X=1195540 $Y=1196130
X2519 11544 25 26 11101 CLKINVX1 $T=1196920 1052470 0 180 $X=1196000 $Y=1048530
X2520 11410 25 26 10427 CLKINVX1 $T=1197380 1229590 1 180 $X=1196460 $Y=1229338
X2521 11135 25 26 11483 CLKINVX1 $T=1196920 1126270 0 0 $X=1196918 $Y=1126018
X2522 10716 25 26 11406 CLKINVX1 $T=1196920 1185310 0 0 $X=1196918 $Y=1185058
X2523 11399 25 26 11420 CLKINVX1 $T=1196920 1340290 0 0 $X=1196918 $Y=1340038
X2524 11262 25 26 11450 CLKINVX1 $T=1198300 1170550 1 0 $X=1198298 $Y=1166610
X2525 10352 25 26 11563 CLKINVX1 $T=1198300 1310770 1 0 $X=1198298 $Y=1306830
X2526 11304 25 26 11451 CLKINVX1 $T=1198300 1310770 0 0 $X=1198298 $Y=1310518
X2527 11965 25 26 11316 CLKINVX1 $T=1199680 1030330 1 180 $X=1198760 $Y=1030078
X2528 11385 25 26 11438 CLKINVX1 $T=1199680 1332910 0 180 $X=1198760 $Y=1328970
X2529 11411 25 26 11454 CLKINVX1 $T=1201060 1325530 0 0 $X=1201058 $Y=1325278
X2530 11463 25 26 11539 CLKINVX1 $T=1203360 1037710 0 0 $X=1203358 $Y=1037458
X2531 11506 25 26 11540 CLKINVX1 $T=1203360 1045090 0 0 $X=1203358 $Y=1044838
X2532 11492 25 26 11542 CLKINVX1 $T=1203360 1303390 1 0 $X=1203358 $Y=1299450
X2533 11505 25 26 11455 CLKINVX1 $T=1204280 1074610 0 180 $X=1203360 $Y=1070670
X2534 10837 25 26 11576 CLKINVX1 $T=1205200 1192690 0 0 $X=1205198 $Y=1192438
X2535 11604 25 26 11419 CLKINVX1 $T=1206120 1318150 1 180 $X=1205200 $Y=1317898
X2536 11175 25 26 11635 CLKINVX1 $T=1205660 1310770 0 0 $X=1205658 $Y=1310518
X2537 11267 25 26 11633 CLKINVX1 $T=1206120 1266490 0 0 $X=1206118 $Y=1266238
X2538 10469 25 26 11556 CLKINVX1 $T=1206580 1096750 0 0 $X=1206578 $Y=1096498
X2539 11686 25 26 11200 CLKINVX1 $T=1208420 1074610 0 180 $X=1207500 $Y=1070670
X2540 11579 25 26 11734 CLKINVX1 $T=1207960 1259110 1 0 $X=1207958 $Y=1255170
X2541 11333 25 26 11625 CLKINVX1 $T=1207960 1318150 1 0 $X=1207958 $Y=1314210
X2542 11311 25 26 11645 CLKINVX1 $T=1208420 1281250 0 0 $X=1208418 $Y=1280998
X2543 11556 25 26 11206 CLKINVX1 $T=1208880 1037710 1 0 $X=1208878 $Y=1033770
X2544 192 25 26 11721 CLKINVX1 $T=1209340 1325530 0 0 $X=1209338 $Y=1325278
X2545 11613 25 26 11582 CLKINVX1 $T=1209800 1067230 1 0 $X=1209798 $Y=1063290
X2546 11522 25 26 11674 CLKINVX1 $T=1209800 1236970 0 0 $X=1209798 $Y=1236718
X2547 11402 25 26 11688 CLKINVX1 $T=1209800 1251730 0 0 $X=1209798 $Y=1251478
X2548 11608 25 26 11659 CLKINVX1 $T=1210720 1081990 0 180 $X=1209800 $Y=1078050
X2549 11575 25 26 11705 CLKINVX1 $T=1210720 1281250 0 0 $X=1210718 $Y=1280998
X2550 10448 25 26 11810 CLKINVX1 $T=1213480 1207450 1 0 $X=1213478 $Y=1203510
X2551 199 25 26 11752 CLKINVX1 $T=1213480 1325530 0 0 $X=1213478 $Y=1325278
X2552 11763 25 26 11488 CLKINVX1 $T=1214860 1037710 0 180 $X=1213940 $Y=1033770
X2553 196 25 26 11729 CLKINVX1 $T=1214860 1281250 1 180 $X=1213940 $Y=1280998
X2554 11437 25 26 11425 CLKINVX1 $T=1214400 1163170 1 0 $X=1214398 $Y=1159230
X2555 9801 25 26 11827 CLKINVX1 $T=1214400 1244350 1 0 $X=1214398 $Y=1240410
X2556 179 25 26 11779 CLKINVX1 $T=1214400 1259110 0 0 $X=1214398 $Y=1258858
X2557 11840 25 26 10480 CLKINVX1 $T=1215320 1200070 1 180 $X=1214400 $Y=1199818
X2558 10107 25 26 11896 CLKINVX1 $T=1215320 1214830 0 0 $X=1215318 $Y=1214578
X2559 9992 25 26 11932 CLKINVX1 $T=1215320 1236970 1 0 $X=1215318 $Y=1233030
X2560 11867 25 26 11879 CLKINVX1 $T=1216240 1037710 1 180 $X=1215320 $Y=1037458
X2561 11323 25 26 11177 CLKINVX1 $T=1215780 1141030 1 0 $X=1215778 $Y=1137090
X2562 11147 25 26 11314 CLKINVX1 $T=1220380 1163170 1 0 $X=1220378 $Y=1159230
X2563 11712 25 26 11894 CLKINVX1 $T=1223140 1052470 0 180 $X=1222220 $Y=1048530
X2564 11322 25 26 11345 CLKINVX1 $T=1223600 1133650 1 0 $X=1223598 $Y=1129710
X2565 206 25 26 11996 CLKINVX1 $T=1224520 1332910 1 0 $X=1224518 $Y=1328970
X2566 11023 25 26 11220 CLKINVX1 $T=1224980 1148410 0 0 $X=1224978 $Y=1148158
X2567 12048 25 26 11529 CLKINVX1 $T=1225900 1052470 1 180 $X=1224980 $Y=1052218
X2568 210 25 26 12010 CLKINVX1 $T=1226820 1332910 0 180 $X=1225900 $Y=1328970
X2569 11786 25 26 11928 CLKINVX1 $T=1226360 1347670 0 0 $X=1226358 $Y=1347418
X2570 12062 25 26 11903 CLKINVX1 $T=1227280 1200070 1 180 $X=1226360 $Y=1199818
X2571 11809 25 26 12131 CLKINVX1 $T=1226820 1096750 1 0 $X=1226818 $Y=1092810
X2572 10967 25 26 11980 CLKINVX1 $T=1227740 1185310 0 0 $X=1227738 $Y=1185058
X2573 12211 25 26 10932 CLKINVX1 $T=1230960 1192690 1 180 $X=1230040 $Y=1192438
X2574 12114 25 26 12106 CLKINVX1 $T=1231420 1236970 1 180 $X=1230500 $Y=1236718
X2575 11868 25 26 12196 CLKINVX1 $T=1230960 1318150 0 0 $X=1230958 $Y=1317898
X2576 11315 25 26 12139 CLKINVX1 $T=1231420 1222210 0 0 $X=1231418 $Y=1221958
X2577 204 25 26 12137 CLKINVX1 $T=1231420 1296010 1 0 $X=1231418 $Y=1292070
X2578 12140 25 26 11860 CLKINVX1 $T=1232340 1067230 0 180 $X=1231420 $Y=1063290
X2579 10533 25 26 12163 CLKINVX1 $T=1232800 1207450 1 0 $X=1232798 $Y=1203510
X2580 10449 25 26 12186 CLKINVX1 $T=1233720 1251730 1 0 $X=1233718 $Y=1247790
X2581 10532 25 26 12193 CLKINVX1 $T=1234180 1192690 1 0 $X=1234178 $Y=1188750
X2582 12219 25 26 12124 CLKINVX1 $T=1236020 1163170 1 180 $X=1235100 $Y=1162918
X2583 216 25 26 12314 CLKINVX1 $T=1236480 1229590 1 0 $X=1236478 $Y=1225650
X2584 10729 25 26 12138 CLKINVX1 $T=1236940 1340290 1 0 $X=1236938 $Y=1336350
X2585 12008 25 26 12077 CLKINVX1 $T=1237400 1170550 0 0 $X=1237398 $Y=1170298
X2586 12256 25 26 12262 CLKINVX1 $T=1237860 1310770 1 0 $X=1237858 $Y=1306830
X2587 12118 25 26 10620 CLKINVX1 $T=1238780 1200070 1 180 $X=1237860 $Y=1199818
X2588 12278 25 26 12231 CLKINVX1 $T=1239700 1118890 0 180 $X=1238780 $Y=1114950
X2589 10670 25 26 12316 CLKINVX1 $T=1240620 1340290 1 0 $X=1240618 $Y=1336350
X2590 12344 25 26 12315 CLKINVX1 $T=1245220 1236970 0 0 $X=1245218 $Y=1236718
X2591 12379 25 26 12404 CLKINVX1 $T=1246140 1192690 1 180 $X=1245220 $Y=1192438
X2592 12297 25 26 12459 CLKINVX1 $T=1245680 1325530 0 0 $X=1245678 $Y=1325278
X2593 12445 25 26 12458 CLKINVX1 $T=1247060 1288630 0 0 $X=1247058 $Y=1288378
X2594 12453 25 26 12460 CLKINVX1 $T=1247980 1067230 0 0 $X=1247978 $Y=1066978
X2595 12454 25 26 12466 CLKINVX1 $T=1247980 1074610 1 0 $X=1247978 $Y=1070670
X2596 12173 25 26 12455 CLKINVX1 $T=1247980 1340290 0 0 $X=1247978 $Y=1340038
X2597 12464 25 26 12449 CLKINVX1 $T=1248900 1059850 0 180 $X=1247980 $Y=1055910
X2598 12303 25 26 12472 CLKINVX1 $T=1248440 1200070 0 0 $X=1248438 $Y=1199818
X2599 12330 25 26 12527 CLKINVX1 $T=1248440 1332910 0 0 $X=1248438 $Y=1332658
X2600 11942 25 26 12366 CLKINVX1 $T=1249360 1303390 0 180 $X=1248440 $Y=1299450
X2601 232 25 26 12506 CLKINVX1 $T=1248900 1347670 1 0 $X=1248898 $Y=1343730
X2602 12503 25 26 11289 CLKINVX1 $T=1249820 1244350 0 180 $X=1248900 $Y=1240410
X2603 12545 25 26 12329 CLKINVX1 $T=1251200 1052470 0 180 $X=1250280 $Y=1048530
X2604 12578 25 26 11162 CLKINVX1 $T=1252120 1200070 0 180 $X=1251200 $Y=1196130
X2605 248 25 26 12634 CLKINVX1 $T=1254420 1347670 1 0 $X=1254418 $Y=1343730
X2606 12604 25 26 12672 CLKINVX1 $T=1254880 1067230 0 0 $X=1254878 $Y=1066978
X2607 12389 25 26 12641 CLKINVX1 $T=1254880 1266490 1 0 $X=1254878 $Y=1262550
X2608 12650 25 26 12600 CLKINVX1 $T=1255800 1067230 0 180 $X=1254880 $Y=1063290
X2609 12642 25 26 12548 CLKINVX1 $T=1255340 1273870 1 0 $X=1255338 $Y=1269930
X2610 12420 25 26 12766 CLKINVX1 $T=1259020 1332910 0 0 $X=1259018 $Y=1332658
X2611 12767 25 26 12701 CLKINVX1 $T=1261320 1200070 1 180 $X=1260400 $Y=1199818
X2612 12829 25 26 12763 CLKINVX1 $T=1261780 1089370 0 180 $X=1260860 $Y=1085430
X2613 12781 25 26 12818 CLKINVX1 $T=1261320 1325530 0 0 $X=1261318 $Y=1325278
X2614 12796 25 26 12780 CLKINVX1 $T=1262240 1185310 0 180 $X=1261320 $Y=1181370
X2615 12706 25 26 12588 CLKINVX1 $T=1262700 1074610 0 180 $X=1261780 $Y=1070670
X2616 12803 25 26 12821 CLKINVX1 $T=1262240 1288630 1 0 $X=1262238 $Y=1284690
X2617 12835 25 26 12912 CLKINVX1 $T=1266380 1340290 0 0 $X=1266378 $Y=1340038
X2618 12881 25 26 12717 CLKINVX1 $T=1267300 1104130 1 180 $X=1266380 $Y=1103878
X2619 12896 25 26 12914 CLKINVX1 $T=1267300 1200070 1 0 $X=1267298 $Y=1196130
X2620 13003 25 26 12716 CLKINVX1 $T=1268680 1081990 1 180 $X=1267760 $Y=1081738
X2621 268 25 26 12964 CLKINVX1 $T=1268220 1347670 0 0 $X=1268218 $Y=1347418
X2622 12232 25 26 12947 CLKINVX1 $T=1268680 1288630 0 0 $X=1268678 $Y=1288378
X2623 276 25 26 11431 CLKINVX1 $T=1270520 1310770 1 180 $X=1269600 $Y=1310518
X2624 12911 25 26 13000 CLKINVX1 $T=1270520 1207450 1 0 $X=1270518 $Y=1203510
X2625 13030 25 26 12849 CLKINVX1 $T=1271440 1104130 0 180 $X=1270520 $Y=1100190
X2626 13054 25 26 12916 CLKINVX1 $T=1273280 1059850 1 180 $X=1272360 $Y=1059598
X2627 13024 25 26 13039 CLKINVX1 $T=1272820 1303390 1 0 $X=1272818 $Y=1299450
X2628 13025 25 26 13098 CLKINVX1 $T=1272820 1310770 1 0 $X=1272818 $Y=1306830
X2629 12694 25 26 13097 CLKINVX1 $T=1273740 1259110 0 0 $X=1273738 $Y=1258858
X2630 12993 25 26 13079 CLKINVX1 $T=1274200 1214830 0 0 $X=1274198 $Y=1214578
X2631 12930 25 26 13118 CLKINVX1 $T=1274200 1222210 1 0 $X=1274198 $Y=1218270
X2632 13008 25 26 13011 CLKINVX1 $T=1275580 1192690 1 0 $X=1275578 $Y=1188750
X2633 283 25 26 13099 CLKINVX1 $T=1277880 1347670 1 180 $X=1276960 $Y=1347418
X2634 12986 25 26 13110 CLKINVX1 $T=1277420 1273870 0 0 $X=1277418 $Y=1273618
X2635 13066 25 26 13129 CLKINVX1 $T=1278800 1244350 1 0 $X=1278798 $Y=1240410
X2636 265 25 26 13238 CLKINVX1 $T=1278800 1259110 0 0 $X=1278798 $Y=1258858
X2637 220 25 26 13220 CLKINVX1 $T=1280640 1332910 0 0 $X=1280638 $Y=1332658
X2638 12945 25 26 13228 CLKINVX1 $T=1281560 1273870 1 0 $X=1281558 $Y=1269930
X2639 13235 25 26 11230 CLKINVX1 $T=1282940 1266490 0 180 $X=1282020 $Y=1262550
X2640 13237 25 26 13159 CLKINVX1 $T=1283400 1185310 1 180 $X=1282480 $Y=1185058
X2641 13183 25 26 13095 CLKINVX1 $T=1282940 1229590 1 0 $X=1282938 $Y=1225650
X2642 13102 25 26 13033 CLKINVX1 $T=1283400 1244350 1 0 $X=1283398 $Y=1240410
X2643 12858 25 26 13258 CLKINVX1 $T=1283400 1266490 1 0 $X=1283398 $Y=1262550
X2644 13251 25 26 13162 CLKINVX1 $T=1284780 1067230 0 180 $X=1283860 $Y=1063290
X2645 13350 25 26 9994 CLKINVX1 $T=1286160 1288630 0 180 $X=1285240 $Y=1284690
X2646 294 25 26 13308 CLKINVX1 $T=1285700 1200070 1 0 $X=1285698 $Y=1196130
X2647 142 25 26 13275 CLKINVX1 $T=1287080 1200070 0 0 $X=1287078 $Y=1199818
X2648 212 25 26 13392 CLKINVX1 $T=1289380 1340290 0 0 $X=1289378 $Y=1340038
X2649 311 25 26 13429 CLKINVX1 $T=1290760 1259110 0 0 $X=1290758 $Y=1258858
X2650 13428 25 26 13385 CLKINVX1 $T=1292600 1148410 1 0 $X=1292598 $Y=1144470
X2651 53 25 26 315 CLKINVX1 $T=1293520 1288630 1 0 $X=1293518 $Y=1284690
X2652 151 25 26 13490 CLKINVX1 $T=1294440 1200070 1 0 $X=1294438 $Y=1196130
X2653 187 25 26 13470 CLKINVX1 $T=1294900 1229590 0 0 $X=1294898 $Y=1229338
X2654 13471 25 26 9922 CLKINVX1 $T=1295820 1296010 0 180 $X=1294900 $Y=1292070
X2655 325 25 26 10792 CLKINVX1 $T=1295820 1310770 0 180 $X=1294900 $Y=1306830
X2656 13448 25 26 13515 CLKINVX1 $T=1296740 1118890 0 0 $X=1296738 $Y=1118638
X2657 326 25 26 13519 CLKINVX1 $T=1296740 1318150 0 0 $X=1296738 $Y=1317898
X2658 291 25 26 13626 CLKINVX1 $T=1297200 1200070 0 0 $X=1297198 $Y=1199818
X2659 13567 25 26 10919 CLKINVX1 $T=1300420 1229590 1 180 $X=1299500 $Y=1229338
X2660 302 25 26 13587 CLKINVX1 $T=1299960 1259110 1 0 $X=1299958 $Y=1255170
X2661 330 25 26 11111 CLKINVX1 $T=1300880 1296010 0 180 $X=1299960 $Y=1292070
X2662 211 25 26 13568 CLKINVX1 $T=1300880 1325530 0 180 $X=1299960 $Y=1321590
X2663 333 25 26 13624 CLKINVX1 $T=1301340 1288630 0 0 $X=1301338 $Y=1288378
X2664 13629 25 26 11202 CLKINVX1 $T=1303180 1296010 0 180 $X=1302260 $Y=1292070
X2665 161 25 26 13639 CLKINVX1 $T=1302720 1200070 0 0 $X=1302718 $Y=1199818
X2666 13506 25 26 13466 CLKINVX1 $T=1303640 1111510 0 180 $X=1302720 $Y=1107570
X2667 13532 25 26 13431 CLKINVX1 $T=1303180 1089370 1 0 $X=1303178 $Y=1085430
X2668 182 25 26 13649 CLKINVX1 $T=1303180 1236970 0 0 $X=1303178 $Y=1236718
X2669 13679 25 26 11114 CLKINVX1 $T=1306400 1288630 1 180 $X=1305480 $Y=1288378
X2670 13562 25 26 13613 CLKINVX1 $T=1306860 1133650 0 0 $X=1306858 $Y=1133398
X2671 13689 25 26 11336 CLKINVX1 $T=1309620 1266490 1 180 $X=1308700 $Y=1266238
X2672 153 25 26 13691 CLKINVX1 $T=1309160 1222210 1 0 $X=1309158 $Y=1218270
X2673 13717 25 26 11285 CLKINVX1 $T=1312380 1273870 1 180 $X=1311460 $Y=1273618
X2674 13418 25 26 13715 CLKINVX1 $T=1311920 1104130 0 0 $X=1311918 $Y=1103878
X2675 13554 25 26 13586 CLKINVX1 $T=1311920 1141030 1 0 $X=1311918 $Y=1137090
X2676 13725 25 26 11374 CLKINVX1 $T=1313300 1266490 0 180 $X=1312380 $Y=1262550
X2677 13739 25 26 11465 CLKINVX1 $T=1314680 1222210 0 180 $X=1313760 $Y=1218270
X2678 13786 25 26 11266 CLKINVX1 $T=1314680 1288630 0 180 $X=1313760 $Y=1284690
X2679 13782 25 26 10296 CLKINVX1 $T=1315140 1207450 1 180 $X=1314220 $Y=1207198
X2680 13764 25 26 10766 CLKINVX1 $T=1316060 1200070 0 180 $X=1315140 $Y=1196130
X2681 355 25 26 10791 CLKINVX1 $T=1320200 1303390 0 180 $X=1319280 $Y=1299450
X2682 13843 25 26 10265 CLKINVX1 $T=1321120 1266490 1 180 $X=1320200 $Y=1266238
X2683 13881 25 26 10095 CLKINVX1 $T=1325720 1222210 0 180 $X=1324800 $Y=1218270
X2684 13902 25 26 11085 CLKINVX1 $T=1327100 1200070 1 180 $X=1326180 $Y=1199818
X2685 13919 25 26 10050 CLKINVX1 $T=1330780 1273870 1 180 $X=1329860 $Y=1273618
X2686 372 25 26 10888 CLKINVX1 $T=1331240 1288630 1 180 $X=1330320 $Y=1288378
X2687 13958 25 26 10626 CLKINVX1 $T=1332160 1200070 1 180 $X=1331240 $Y=1199818
X2688 13971 25 26 10588 CLKINVX1 $T=1334920 1273870 0 180 $X=1334000 $Y=1269930
X2689 395 25 26 11216 CLKINVX1 $T=1339520 1310770 0 180 $X=1338600 $Y=1306830
X2690 14203 25 26 10074 CLKINVX1 $T=1354240 1236970 1 180 $X=1353320 $Y=1236718
X2691 14458 25 26 10571 CLKINVX1 $T=1373100 1214830 0 180 $X=1372180 $Y=1210890
X2692 14741 25 26 11310 CLKINVX1 $T=1402080 1296010 0 180 $X=1401160 $Y=1292070
X2693 14743 25 26 10454 CLKINVX1 $T=1402540 1251730 0 180 $X=1401620 $Y=1247790
X2694 14833 25 26 10402 CLKINVX1 $T=1411740 1200070 1 180 $X=1410820 $Y=1199818
X2695 13726 25 26 625 CLKINVX1 $T=1608620 1332910 0 0 $X=1608618 $Y=1332658
X2696 13726 25 26 619 CLKINVX1 $T=1614140 1340290 1 0 $X=1614138 $Y=1336350
X2697 8945 26 25 8919 INVXL $T=1063060 1104130 1 180 $X=1062140 $Y=1103878
X2698 8903 26 25 8973 INVXL $T=1064900 1081990 0 0 $X=1064898 $Y=1081738
X2699 8864 26 25 9041 INVXL $T=1069960 1185310 0 0 $X=1069958 $Y=1185058
X2700 9014 26 25 9037 INVXL $T=1070880 1089370 1 0 $X=1070878 $Y=1085430
X2701 8871 26 25 9006 INVXL $T=1070880 1192690 0 0 $X=1070878 $Y=1192438
X2702 9085 26 25 9073 INVXL $T=1075940 1111510 0 180 $X=1075020 $Y=1107570
X2703 9008 26 25 9002 INVXL $T=1078700 1074610 1 180 $X=1077780 $Y=1074358
X2704 9105 26 25 9312 INVXL $T=1081460 1052470 0 0 $X=1081458 $Y=1052218
X2705 9078 26 25 9242 INVXL $T=1081920 1133650 1 0 $X=1081918 $Y=1129710
X2706 9118 26 25 9245 INVXL $T=1082380 1096750 0 0 $X=1082378 $Y=1096498
X2707 9153 26 25 9227 INVXL $T=1082380 1104130 1 0 $X=1082378 $Y=1100190
X2708 9271 26 25 9257 INVXL $T=1088360 1141030 1 180 $X=1087440 $Y=1140778
X2709 9355 26 25 9439 INVXL $T=1094340 1096750 1 0 $X=1094338 $Y=1092810
X2710 9405 26 25 9381 INVXL $T=1096180 1318150 1 180 $X=1095260 $Y=1317898
X2711 9362 26 25 9389 INVXL $T=1098020 1104130 1 180 $X=1097100 $Y=1103878
X2712 46 26 25 9663 INVXL $T=1098020 1288630 1 0 $X=1098018 $Y=1284690
X2713 9217 26 25 9467 INVXL $T=1100320 1133650 1 0 $X=1100318 $Y=1129710
X2714 9415 26 25 9506 INVXL $T=1100780 1148410 1 0 $X=1100778 $Y=1144470
X2715 9475 26 25 9597 INVXL $T=1101700 1074610 0 0 $X=1101698 $Y=1074358
X2716 9381 26 25 57 INVXL $T=1104000 1318150 0 0 $X=1103998 $Y=1317898
X2717 9151 26 25 9428 INVXL $T=1106300 1229590 0 0 $X=1106298 $Y=1229338
X2718 9283 26 25 9259 INVXL $T=1109520 1200070 0 0 $X=1109518 $Y=1199818
X2719 9097 26 25 9680 INVXL $T=1109980 1192690 0 0 $X=1109978 $Y=1192438
X2720 57 26 25 9558 INVXL $T=1109980 1340290 1 0 $X=1109978 $Y=1336350
X2721 9138 26 25 9779 INVXL $T=1110440 1118890 0 0 $X=1110438 $Y=1118638
X2722 8885 26 25 9678 INVXL $T=1110440 1141030 1 0 $X=1110438 $Y=1137090
X2723 9785 26 25 9824 INVXL $T=1115040 1089370 0 0 $X=1115038 $Y=1089118
X2724 9061 26 25 9836 INVXL $T=1116420 1155790 1 0 $X=1116418 $Y=1151850
X2725 8834 26 25 9812 INVXL $T=1116880 1163170 0 0 $X=1116878 $Y=1162918
X2726 9238 26 25 9884 INVXL $T=1122860 1126270 0 180 $X=1121940 $Y=1122330
X2727 9714 26 25 9869 INVXL $T=1123780 1045090 0 180 $X=1122860 $Y=1041150
X2728 79 26 25 9929 INVXL $T=1123320 1318150 1 0 $X=1123318 $Y=1314210
X2729 88 26 25 9953 INVXL $T=1127460 1318150 0 0 $X=1127458 $Y=1317898
X2730 9893 26 25 10016 INVXL $T=1129300 1045090 0 180 $X=1128380 $Y=1041150
X2731 8917 26 25 10057 INVXL $T=1129300 1141030 1 180 $X=1128380 $Y=1140778
X2732 8964 26 25 10061 INVXL $T=1130680 1155790 1 180 $X=1129760 $Y=1155538
X2733 9258 26 25 10211 INVXL $T=1134360 1126270 0 0 $X=1134358 $Y=1126018
X2734 9534 26 25 10412 INVXL $T=1144940 1155790 1 0 $X=1144938 $Y=1151850
X2735 9512 26 25 10332 INVXL $T=1146320 1148410 0 180 $X=1145400 $Y=1144470
X2736 9806 26 25 9918 INVXL $T=1151840 1141030 0 0 $X=1151838 $Y=1140778
X2737 10136 26 25 9952 INVXL $T=1154600 1185310 1 0 $X=1154598 $Y=1181370
X2738 9386 26 25 10435 INVXL $T=1157360 1148410 1 0 $X=1157358 $Y=1144470
X2739 10740 26 25 10675 INVXL $T=1162420 1096750 0 180 $X=1161500 $Y=1092810
X2740 9270 26 25 10602 INVXL $T=1163340 1126270 1 180 $X=1162420 $Y=1126018
X2741 10583 26 25 10865 INVXL $T=1167940 1045090 1 0 $X=1167938 $Y=1041150
X2742 10920 26 25 148 INVXL $T=1172540 1347670 0 0 $X=1172538 $Y=1347418
X2743 10995 26 25 11076 INVXL $T=1178520 1170550 1 0 $X=1178518 $Y=1166610
X2744 11254 26 25 11273 INVXL $T=1188180 1347670 1 0 $X=1188178 $Y=1343730
X2745 11149 26 25 11245 INVXL $T=1188640 1325530 1 0 $X=1188638 $Y=1321590
X2746 11380 26 25 10669 INVXL $T=1191860 1281250 0 180 $X=1190940 $Y=1277310
X2747 11355 26 25 11380 INVXL $T=1194160 1273870 0 0 $X=1194158 $Y=1273618
X2748 11391 26 25 11399 INVXL $T=1196920 1340290 0 180 $X=1196000 $Y=1336350
X2749 11422 26 25 11605 INVXL $T=1205200 1325530 0 0 $X=1205198 $Y=1325278
X2750 10967 26 25 11449 INVXL $T=1208880 1148410 0 0 $X=1208878 $Y=1148158
X2751 11546 26 25 11591 INVXL $T=1209800 1185310 1 180 $X=1208880 $Y=1185058
X2752 11764 26 25 11616 INVXL $T=1210720 1096750 1 180 $X=1209800 $Y=1096498
X2753 11749 26 25 11740 INVXL $T=1214400 1111510 0 180 $X=1213480 $Y=1107570
X2754 11052 26 25 11561 INVXL $T=1216240 1185310 0 0 $X=1216238 $Y=1185058
X2755 111 26 25 11891 INVXL $T=1216700 1207450 1 0 $X=1216698 $Y=1203510
X2756 109 26 25 11991 INVXL $T=1219920 1303390 0 0 $X=1219918 $Y=1303138
X2757 11732 26 25 11816 INVXL $T=1220840 1104130 1 180 $X=1219920 $Y=1103878
X2758 70 26 25 11977 INVXL $T=1220840 1288630 1 0 $X=1220838 $Y=1284690
X2759 40 26 25 11978 INVXL $T=1220840 1318150 1 0 $X=1220838 $Y=1314210
X2760 11798 26 25 11817 INVXL $T=1224980 1118890 0 0 $X=1224978 $Y=1118638
X2761 11984 26 25 11818 INVXL $T=1224980 1185310 1 0 $X=1224978 $Y=1181370
X2762 51 26 25 12009 INVXL $T=1225440 1273870 1 0 $X=1225438 $Y=1269930
X2763 11926 26 25 12013 INVXL $T=1226360 1163170 1 0 $X=1226358 $Y=1159230
X2764 11901 26 25 11874 INVXL $T=1227740 1133650 1 180 $X=1226820 $Y=1133398
X2765 87 26 25 11988 INVXL $T=1227740 1244350 0 180 $X=1226820 $Y=1240410
X2766 75 26 25 11990 INVXL $T=1227740 1259110 1 180 $X=1226820 $Y=1258858
X2767 80 26 25 11989 INVXL $T=1230960 1251730 0 180 $X=1230040 $Y=1247790
X2768 12116 26 25 11324 INVXL $T=1230960 1288630 0 180 $X=1230040 $Y=1284690
X2769 11941 26 25 11828 INVXL $T=1230500 1170550 0 0 $X=1230498 $Y=1170298
X2770 12125 26 25 11060 INVXL $T=1231880 1273870 1 180 $X=1230960 $Y=1273618
X2771 55 26 25 12119 INVXL $T=1231420 1229590 1 0 $X=1231418 $Y=1225650
X2772 11821 26 25 12116 INVXL $T=1233260 1281250 0 180 $X=1232340 $Y=1277310
X2773 100 26 25 12038 INVXL $T=1232800 1222210 1 0 $X=1232798 $Y=1218270
X2774 12236 26 25 12157 INVXL $T=1234180 1111510 1 180 $X=1233260 $Y=1111258
X2775 45 26 25 12260 INVXL $T=1235100 1296010 0 0 $X=1235098 $Y=1295758
X2776 12223 26 25 12121 INVXL $T=1236020 1104130 0 180 $X=1235100 $Y=1100190
X2777 12154 26 25 12214 INVXL $T=1236020 1141030 1 180 $X=1235100 $Y=1140778
X2778 12259 26 25 12125 INVXL $T=1236020 1273870 1 180 $X=1235100 $Y=1273618
X2779 12251 26 25 11025 INVXL $T=1237400 1259110 1 0 $X=1237398 $Y=1255170
X2780 12221 26 25 12251 INVXL $T=1238320 1251730 1 180 $X=1237400 $Y=1251478
X2781 12253 26 25 12191 INVXL $T=1238780 1133650 1 0 $X=1238778 $Y=1129710
X2782 139 26 25 12323 INVXL $T=1240620 1207450 1 0 $X=1240618 $Y=1203510
X2783 12266 26 25 12267 INVXL $T=1243380 1118890 1 180 $X=1242460 $Y=1118638
X2784 56 26 25 12171 INVXL $T=1243380 1266490 1 180 $X=1242460 $Y=1266238
X2785 12393 26 25 12285 INVXL $T=1244760 1133650 1 180 $X=1243840 $Y=1133398
X2786 177 26 25 12284 INVXL $T=1245220 1318150 1 180 $X=1244300 $Y=1317898
X2787 12498 26 25 11228 INVXL $T=1248900 1273870 1 180 $X=1247980 $Y=1273618
X2788 12333 26 25 12367 INVXL $T=1249360 1104130 1 180 $X=1248440 $Y=1103878
X2789 12249 26 25 12382 INVXL $T=1249360 1163170 0 180 $X=1248440 $Y=1159230
X2790 11728 26 25 12514 INVXL $T=1248900 1177930 1 0 $X=1248898 $Y=1173990
X2791 12405 26 25 12498 INVXL $T=1248900 1266490 1 0 $X=1248898 $Y=1262550
X2792 12529 26 25 10969 INVXL $T=1250280 1281250 1 0 $X=1250278 $Y=1277310
X2793 12581 26 25 12529 INVXL $T=1251200 1273870 1 180 $X=1250280 $Y=1273618
X2794 12596 26 25 12578 INVXL $T=1253500 1200070 1 180 $X=1252580 $Y=1199818
X2795 231 26 25 12617 INVXL $T=1254880 1332910 1 0 $X=1254878 $Y=1328970
X2796 12691 26 25 12631 INVXL $T=1255800 1089370 0 180 $X=1254880 $Y=1085430
X2797 117 26 25 12599 INVXL $T=1255800 1244350 0 180 $X=1254880 $Y=1240410
X2798 12702 26 25 10987 INVXL $T=1257180 1244350 1 180 $X=1256260 $Y=1244098
X2799 12704 26 25 12722 INVXL $T=1258560 1045090 0 0 $X=1258558 $Y=1044838
X2800 11275 26 25 12463 INVXL $T=1260860 1118890 0 0 $X=1260858 $Y=1118638
X2801 213 26 25 12727 INVXL $T=1261780 1303390 1 180 $X=1260860 $Y=1303138
X2802 12795 26 25 11108 INVXL $T=1262240 1200070 1 180 $X=1261320 $Y=1199818
X2803 124 26 25 12649 INVXL $T=1262240 1214830 0 180 $X=1261320 $Y=1210890
X2804 143 26 25 12726 INVXL $T=1262700 1222210 0 180 $X=1261780 $Y=1218270
X2805 12500 26 25 12678 INVXL $T=1263160 1148410 0 180 $X=1262240 $Y=1144470
X2806 12843 26 25 11416 INVXL $T=1264540 1192690 1 180 $X=1263620 $Y=1192438
X2807 12844 26 25 11229 INVXL $T=1264540 1214830 0 180 $X=1263620 $Y=1210890
X2808 12866 26 25 11186 INVXL $T=1265460 1185310 1 180 $X=1264540 $Y=1185058
X2809 12876 26 25 12843 INVXL $T=1265460 1192690 1 180 $X=1264540 $Y=1192438
X2810 12877 26 25 12844 INVXL $T=1265460 1214830 0 180 $X=1264540 $Y=1210890
X2811 12867 26 25 12795 INVXL $T=1265920 1200070 0 180 $X=1265000 $Y=1196130
X2812 11244 26 25 12622 INVXL $T=1265920 1133650 1 0 $X=1265918 $Y=1129710
X2813 12582 26 25 12863 INVXL $T=1266840 1170550 1 180 $X=1265920 $Y=1170298
X2814 12878 26 25 10986 INVXL $T=1266840 1222210 0 180 $X=1265920 $Y=1218270
X2815 12762 26 25 12869 INVXL $T=1267300 1067230 0 180 $X=1266380 $Y=1063290
X2816 12880 26 25 12870 INVXL $T=1267300 1089370 1 180 $X=1266380 $Y=1089118
X2817 12892 26 25 11188 INVXL $T=1267300 1244350 0 180 $X=1266380 $Y=1240410
X2818 12685 26 25 12965 INVXL $T=1267300 1148410 0 0 $X=1267298 $Y=1148158
X2819 13032 26 25 12878 INVXL $T=1268220 1214830 1 180 $X=1267300 $Y=1214578
X2820 12962 26 25 12892 INVXL $T=1268220 1236970 1 180 $X=1267300 $Y=1236718
X2821 13043 26 25 12702 INVXL $T=1270980 1222210 0 180 $X=1270060 $Y=1218270
X2822 227 26 25 12728 INVXL $T=1272820 1318150 1 180 $X=1271900 $Y=1317898
X2823 13056 26 25 12866 INVXL $T=1275120 1177930 1 180 $X=1274200 $Y=1177678
X2824 11066 26 25 12889 INVXL $T=1276500 1141030 1 0 $X=1276498 $Y=1137090
X2825 235 26 25 13119 INVXL $T=1277420 1332910 1 0 $X=1277418 $Y=1328970
X2826 11344 26 25 12874 INVXL $T=1278340 1141030 0 0 $X=1278338 $Y=1140778
X2827 13104 26 25 13107 INVXL $T=1279720 1052470 0 180 $X=1278800 $Y=1048530
X2828 13058 26 25 13147 INVXL $T=1279260 1104130 1 0 $X=1279258 $Y=1100190
X2829 12814 26 25 13065 INVXL $T=1282480 1170550 0 180 $X=1281560 $Y=1166610
X2830 12943 26 25 13055 INVXL $T=1282940 1163170 1 180 $X=1282020 $Y=1162918
X2831 11063 26 25 13346 INVXL $T=1283400 1155790 0 0 $X=1283398 $Y=1155538
X2832 264 26 25 13120 INVXL $T=1284320 1340290 0 180 $X=1283400 $Y=1336350
X2833 11063 26 25 13161 INVXL $T=1283860 1059850 1 0 $X=1283858 $Y=1055910
X2834 11225 26 25 12926 INVXL $T=1284320 1111510 1 0 $X=1284318 $Y=1107570
X2835 241 26 25 13160 INVXL $T=1285240 1318150 0 180 $X=1284320 $Y=1314210
X2836 11087 26 25 12744 INVXL $T=1284780 1111510 0 0 $X=1284778 $Y=1111258
X2837 300 26 25 13295 INVXL $T=1285240 1273870 0 0 $X=1285238 $Y=1273618
X2838 11295 26 25 12729 INVXL $T=1285700 1148410 0 0 $X=1285698 $Y=1148158
X2839 284 26 25 13239 INVXL $T=1285700 1303390 0 0 $X=1285698 $Y=1303138
X2840 13297 26 25 13047 INVXL $T=1286620 1052470 1 180 $X=1285700 $Y=1052218
X2841 289 26 25 13294 INVXL $T=1286160 1236970 0 0 $X=1286158 $Y=1236718
X2842 13389 26 25 13246 INVXL $T=1287540 1089370 1 180 $X=1286620 $Y=1089118
X2843 11243 26 25 12927 INVXL $T=1288460 1126270 1 0 $X=1288458 $Y=1122330
X2844 309 26 25 13296 INVXL $T=1289380 1296010 1 180 $X=1288460 $Y=1295758
X2845 12730 26 25 12941 INVXL $T=1289380 1133650 1 0 $X=1289378 $Y=1129710
X2846 12857 26 25 12955 INVXL $T=1289840 1126270 0 0 $X=1289838 $Y=1126018
X2847 13307 26 25 13463 INVXL $T=1290300 1074610 0 0 $X=1290298 $Y=1074358
X2848 11421 26 25 13453 INVXL $T=1290300 1111510 1 0 $X=1290298 $Y=1107570
X2849 12834 26 25 12815 INVXL $T=1290300 1163170 1 0 $X=1290298 $Y=1159230
X2850 242 26 25 13245 INVXL $T=1291220 1325530 0 180 $X=1290300 $Y=1321590
X2851 279 26 25 13292 INVXL $T=1292140 1229590 0 180 $X=1291220 $Y=1225650
X2852 12929 26 25 13010 INVXL $T=1295360 1148410 1 180 $X=1294440 $Y=1148158
X2853 308 26 25 13305 INVXL $T=1295820 1259110 0 180 $X=1294900 $Y=1255170
X2854 280 26 25 13306 INVXL $T=1295820 1288630 1 180 $X=1294900 $Y=1288378
X2855 13236 26 25 13499 INVXL $T=1296280 1059850 1 0 $X=1296278 $Y=1055910
X2856 13501 26 25 13494 INVXL $T=1297200 1141030 0 180 $X=1296280 $Y=1137090
X2857 13372 26 25 13454 INVXL $T=1297200 1089370 0 0 $X=1297198 $Y=1089118
X2858 12700 26 25 13516 INVXL $T=1302260 1133650 1 0 $X=1302258 $Y=1129710
X2859 13362 26 25 13708 INVXL $T=1303180 1104130 0 0 $X=1303178 $Y=1103878
X2860 321 26 25 13282 INVXL $T=1304560 1266490 1 180 $X=1303640 $Y=1266238
X2861 13261 26 25 13473 INVXL $T=1309160 1074610 1 0 $X=1309158 $Y=1070670
X2862 13393 26 25 13711 INVXL $T=1311920 1081990 0 0 $X=1311918 $Y=1081738
X2863 13582 26 25 13705 INVXL $T=1314220 1111510 0 0 $X=1314218 $Y=1111258
X2864 15981 26 25 16048 INVXL $T=1532720 1148410 1 0 $X=1532718 $Y=1144470
X2865 8748 25 26 8827 INVX1 $T=1052480 1141030 1 0 $X=1052478 $Y=1137090
X2866 8814 25 26 8870 INVX1 $T=1058920 1141030 1 0 $X=1058918 $Y=1137090
X2867 8816 25 26 8931 INVX1 $T=1060300 1133650 1 0 $X=1060298 $Y=1129710
X2868 8961 25 26 9005 INVX1 $T=1082840 1111510 0 0 $X=1082838 $Y=1111258
X2869 9003 25 26 8980 INVX1 $T=1088360 1111510 0 0 $X=1088358 $Y=1111258
X2870 9101 25 26 9243 INVX1 $T=1104000 1133650 0 0 $X=1103998 $Y=1133398
X2871 9509 25 26 9170 INVX1 $T=1130220 1207450 0 180 $X=1129300 $Y=1203510
X2872 9102 25 26 9518 INVX1 $T=1138500 1155790 0 0 $X=1138498 $Y=1155538
X2873 9228 25 26 9437 INVX1 $T=1146320 1133650 1 180 $X=1145400 $Y=1133398
X2874 10530 25 26 10469 INVX1 $T=1155980 1177930 1 0 $X=1155978 $Y=1173990
X2875 10616 25 26 10605 INVX1 $T=1160580 1170550 0 0 $X=1160578 $Y=1170298
X2876 10803 25 26 10877 INVX1 $T=1170700 1170550 0 180 $X=1169780 $Y=1166610
X2877 10595 25 26 10619 INVX1 $T=1174840 1170550 1 0 $X=1174838 $Y=1166610
X2878 10634 25 26 11051 INVX1 $T=1175300 1118890 1 0 $X=1175298 $Y=1114950
X2879 162 25 26 11103 INVX1 $T=1184960 1318150 1 180 $X=1184040 $Y=1317898
X2880 11312 25 26 11122 INVX1 $T=1188640 1318150 1 180 $X=1187720 $Y=1317898
X2881 11397 25 26 11297 INVX1 $T=1194160 1347670 1 180 $X=1193240 $Y=1347418
X2882 11484 25 26 11187 INVX1 $T=1198760 1251730 0 180 $X=1197840 $Y=1247790
X2883 11398 25 26 11725 INVX1 $T=1211180 1074610 1 0 $X=1211178 $Y=1070670
X2884 189 25 26 11756 INVX1 $T=1213940 1259110 1 0 $X=1213938 $Y=1255170
X2885 11773 25 26 11647 INVX1 $T=1215320 1303390 1 180 $X=1214400 $Y=1303138
X2886 11782 25 26 11802 INVX1 $T=1215320 1207450 0 0 $X=1215318 $Y=1207198
X2887 11783 25 26 11803 INVX1 $T=1215320 1229590 0 0 $X=1215318 $Y=1229338
X2888 208 25 26 11210 INVX1 $T=1218080 1340290 1 180 $X=1217160 $Y=1340038
X2889 11871 25 26 11919 INVX1 $T=1219460 1222210 1 0 $X=1219458 $Y=1218270
X2890 11819 25 26 11918 INVX1 $T=1220380 1200070 0 0 $X=1220378 $Y=1199818
X2891 11831 25 26 11893 INVX1 $T=1220840 1244350 0 0 $X=1220838 $Y=1244098
X2892 11929 25 26 11820 INVX1 $T=1221760 1214830 0 180 $X=1220840 $Y=1210890
X2893 11960 25 26 11841 INVX1 $T=1223600 1222210 0 180 $X=1222680 $Y=1218270
X2894 12135 25 26 11291 INVX1 $T=1230960 1259110 1 180 $X=1230040 $Y=1258858
X2895 12215 25 26 11222 INVX1 $T=1232340 1244350 0 180 $X=1231420 $Y=1240410
X2896 12238 25 26 11318 INVX1 $T=1232800 1251730 1 180 $X=1231880 $Y=1251478
X2897 12195 25 26 11292 INVX1 $T=1232800 1259110 0 180 $X=1231880 $Y=1255170
X2898 11993 25 26 12240 INVX1 $T=1234640 1318150 0 0 $X=1234638 $Y=1317898
X2899 12220 25 26 12245 INVX1 $T=1236480 1244350 1 0 $X=1236478 $Y=1240410
X2900 217 25 26 11967 INVX1 $T=1237400 1296010 0 180 $X=1236480 $Y=1292070
X2901 12335 25 26 11427 INVX1 $T=1242460 1229590 0 180 $X=1241540 $Y=1225650
X2902 12224 25 26 12305 INVX1 $T=1242460 1214830 1 0 $X=1242458 $Y=1210890
X2903 12580 25 26 10933 INVX1 $T=1249360 1236970 1 180 $X=1248440 $Y=1236718
X2904 12381 25 26 12546 INVX1 $T=1248900 1089370 1 0 $X=1248898 $Y=1085430
X2905 12473 25 26 12504 INVX1 $T=1248900 1303390 0 0 $X=1248898 $Y=1303138
X2906 12505 25 26 12519 INVX1 $T=1249360 1325530 0 0 $X=1249358 $Y=1325278
X2907 12555 25 26 12562 INVX1 $T=1251200 1340290 0 0 $X=1251198 $Y=1340038
X2908 12565 25 26 11136 INVX1 $T=1253040 1192690 1 180 $X=1252120 $Y=1192438
X2909 12626 25 26 11163 INVX1 $T=1254880 1288630 0 180 $X=1253960 $Y=1284690
X2910 12718 25 26 12607 INVX1 $T=1255800 1303390 1 180 $X=1254880 $Y=1303138
X2911 236 25 26 12856 INVX1 $T=1260860 1244350 1 0 $X=1260858 $Y=1240410
X2912 12819 25 26 12883 INVX1 $T=1266380 1340290 1 0 $X=1266378 $Y=1336350
X2913 12985 25 26 13016 INVX1 $T=1271440 1273870 1 0 $X=1271438 $Y=1269930
X2914 13005 25 26 13046 INVX1 $T=1271440 1340290 0 0 $X=1271438 $Y=1340038
X2915 13057 25 26 12995 INVX1 $T=1272360 1332910 1 180 $X=1271440 $Y=1332658
X2916 12963 25 26 13038 INVX1 $T=1272820 1229590 1 0 $X=1272818 $Y=1225650
X2917 13249 25 26 12957 INVX1 $T=1283860 1273870 0 180 $X=1282940 $Y=1269930
X2918 13264 25 26 12793 INVX1 $T=1284780 1340290 1 180 $X=1283860 $Y=1340038
X2919 13284 25 26 12944 INVX1 $T=1288000 1229590 0 180 $X=1287080 $Y=1225650
X2920 327 25 26 11737 INVX1 $T=1298120 1347670 1 180 $X=1297200 $Y=1347418
X2921 13595 25 26 13718 INVX1 $T=1301800 1081990 0 180 $X=1300880 $Y=1078050
X2922 13628 25 26 10248 INVX1 $T=1303180 1281250 1 180 $X=1302260 $Y=1280998
X2923 13588 25 26 13714 INVX1 $T=1307320 1096750 1 0 $X=1307318 $Y=1092810
X2924 327 25 26 12452 INVX1 $T=1307320 1288630 1 0 $X=1307318 $Y=1284690
X2925 13718 25 26 13367 INVX1 $T=1312840 1067230 1 180 $X=1311920 $Y=1066978
X2926 13811 25 26 10546 INVX1 $T=1318820 1288630 0 180 $X=1317900 $Y=1284690
X2927 14698 25 26 14518 INVX1 $T=1397940 1200070 0 0 $X=1397938 $Y=1199818
X2928 14837 25 26 14698 INVX1 $T=1411740 1200070 0 0 $X=1411738 $Y=1199818
X2929 398 25 26 16121 INVX1 $T=1544220 1148410 1 180 $X=1543300 $Y=1148158
X2930 9329 25 27 26 CLKINVX3 $T=1092960 1251730 1 0 $X=1092958 $Y=1247790
X2931 9316 25 38 26 CLKINVX3 $T=1093880 1207450 0 0 $X=1093878 $Y=1207198
X2932 9549 25 47 26 CLKINVX3 $T=1100780 1207450 1 180 $X=1099400 $Y=1207198
X2933 9488 25 58 26 CLKINVX3 $T=1105380 1214830 1 0 $X=1105378 $Y=1210890
X2934 9651 25 63 26 CLKINVX3 $T=1109520 1214830 1 0 $X=1109518 $Y=1210890
X2935 102 25 10907 26 CLKINVX3 $T=1167940 1340290 0 0 $X=1167938 $Y=1340038
X2936 13350 25 230 26 CLKINVX3 $T=1287540 1296010 1 180 $X=1286160 $Y=1295758
X2937 329 25 13684 26 CLKINVX3 $T=1299960 1340290 0 0 $X=1299958 $Y=1340038
X2938 13628 25 12051 26 CLKINVX3 $T=1316060 1288630 0 0 $X=1316058 $Y=1288378
X2939 379 25 14007 26 CLKINVX3 $T=1331240 1347670 1 0 $X=1331238 $Y=1343730
X2940 53 25 408 26 CLKINVX3 $T=1352860 1192690 1 0 $X=1352858 $Y=1188750
X2941 440 25 441 26 CLKINVX3 $T=1375400 1170550 1 0 $X=1375398 $Y=1166610
X2942 13782 25 12142 26 CLKINVX3 $T=1378160 1214830 0 0 $X=1378158 $Y=1214578
X2943 13471 25 218 26 CLKINVX3 $T=1383680 1318150 1 0 $X=1383678 $Y=1314210
X2944 13811 25 12024 26 CLKINVX3 $T=1384600 1310770 1 0 $X=1384598 $Y=1306830
X2945 456 25 457 26 CLKINVX3 $T=1391960 1170550 0 0 $X=1391958 $Y=1170298
X2946 461 25 464 26 CLKINVX3 $T=1403460 1141030 1 0 $X=1403458 $Y=1137090
X2947 13786 25 317 26 CLKINVX3 $T=1404380 1303390 0 0 $X=1404378 $Y=1303138
X2948 14203 25 12143 26 CLKINVX3 $T=1405760 1229590 0 0 $X=1405758 $Y=1229338
X2949 13629 25 287 26 CLKINVX3 $T=1406680 1347670 1 0 $X=1406678 $Y=1343730
X2950 13881 25 12039 26 CLKINVX3 $T=1416800 1236970 1 0 $X=1416798 $Y=1233030
X2951 13902 25 12792 26 CLKINVX3 $T=1417720 1207450 0 0 $X=1417718 $Y=1207198
X2952 395 25 305 26 CLKINVX3 $T=1419100 1347670 1 0 $X=1419098 $Y=1343730
X2953 325 25 260 26 CLKINVX3 $T=1420480 1325530 1 0 $X=1420478 $Y=1321590
X2954 372 25 228 26 CLKINVX3 $T=1420480 1325530 0 0 $X=1420478 $Y=1325278
X2955 14833 25 12063 26 CLKINVX3 $T=1420940 1207450 0 0 $X=1420938 $Y=1207198
X2956 330 25 252 26 CLKINVX3 $T=1421860 1347670 0 0 $X=1421858 $Y=1347418
X2957 13679 25 296 26 CLKINVX3 $T=1422780 1325530 0 0 $X=1422778 $Y=1325278
X2958 14743 25 12050 26 CLKINVX3 $T=1423240 1251730 1 0 $X=1423238 $Y=1247790
X2959 276 25 262 26 CLKINVX3 $T=1423240 1332910 1 0 $X=1423238 $Y=1328970
X2960 13958 25 12754 26 CLKINVX3 $T=1426920 1207450 1 0 $X=1426918 $Y=1203510
X2961 13971 25 219 26 CLKINVX3 $T=1428760 1273870 1 0 $X=1428758 $Y=1269930
X2962 13919 25 12110 26 CLKINVX3 $T=1433820 1288630 0 0 $X=1433818 $Y=1288378
X2963 355 25 285 26 CLKINVX3 $T=1434280 1347670 0 0 $X=1434278 $Y=1347418
X2964 14741 25 313 26 CLKINVX3 $T=1434740 1303390 1 0 $X=1434738 $Y=1299450
X2965 13764 25 12516 26 CLKINVX3 $T=1436120 1214830 1 0 $X=1436118 $Y=1210890
X2966 14458 25 12589 26 CLKINVX3 $T=1436580 1236970 0 0 $X=1436578 $Y=1236718
X2967 13689 25 13390 26 CLKINVX3 $T=1438880 1266490 0 0 $X=1438878 $Y=1266238
X2968 13843 25 12258 26 CLKINVX3 $T=1438880 1273870 1 0 $X=1438878 $Y=1269930
X2969 13567 25 13405 26 CLKINVX3 $T=1439800 1229590 1 0 $X=1439798 $Y=1225650
X2970 13235 25 299 26 CLKINVX3 $T=1439800 1318150 0 0 $X=1439798 $Y=1317898
X2971 13725 25 13329 26 CLKINVX3 $T=1442560 1266490 0 0 $X=1442558 $Y=1266238
X2972 13717 25 307 26 CLKINVX3 $T=1451760 1310770 1 0 $X=1451758 $Y=1306830
X2973 13739 25 13332 26 CLKINVX3 $T=1456820 1222210 0 0 $X=1456818 $Y=1221958
X2974 16095 25 576 26 CLKINVX3 $T=1566300 1310770 1 0 $X=1566298 $Y=1306830
X2975 492 25 15158 26 CLKBUFX20 $T=1435200 1229590 0 0 $X=1435198 $Y=1229338
X2976 492 25 13676 26 CLKBUFX20 $T=1455440 1318150 1 0 $X=1455438 $Y=1314210
X2977 492 25 15374 26 CLKBUFX20 $T=1455900 1244350 1 0 $X=1455898 $Y=1240410
X2978 26 332 12051 13611 13618 25 13081 13618 13612 12746 306 13518 13591 13740 3920 ICV_28 $T=1299500 1310770 1 0 $X=1299498 $Y=1306830
X2979 26 335 13405 13678 13685 25 13349 13491 13652 11826 306 13744 13623 13816 3920 ICV_28 $T=1304560 1229590 1 0 $X=1304558 $Y=1225650
X2980 26 335 12792 13768 13803 25 13560 13803 13817 11826 338 13354 13815 13988 3920 ICV_28 $T=1315140 1177930 0 0 $X=1315138 $Y=1177678
X2981 26 347 12792 13800 13808 25 13640 13801 13800 13599 342 13906 13808 13954 3920 ICV_28 $T=1315600 1126270 1 0 $X=1315598 $Y=1122330
X2982 26 319 13405 13810 13742 25 13609 13867 13873 13687 339 13744 13856 13965 3920 ICV_28 $T=1319740 1229590 1 0 $X=1319738 $Y=1225650
X2983 26 384 12110 13964 13985 25 13566 14005 13964 12746 362 13736 13985 14108 3920 ICV_28 $T=1332620 1288630 0 0 $X=1332618 $Y=1288378
X2984 26 358 12258 14021 14038 25 348 13922 14021 396 397 13890 14038 14139 3920 ICV_28 $T=1335840 1340290 0 0 $X=1335838 $Y=1340038
X2985 26 347 12142 14040 14047 25 13640 14047 14026 13599 339 13906 14027 14147 3920 ICV_28 $T=1336760 1126270 1 0 $X=1336758 $Y=1122330
X2986 26 350 13332 14057 14042 25 13609 14085 14057 13687 13851 13744 14042 14187 3920 ICV_28 $T=1337680 1222210 0 0 $X=1337678 $Y=1221958
X2987 26 384 230 14086 14032 25 348 14038 14086 396 362 13890 14032 403 3920 ICV_28 $T=1339060 1347670 1 0 $X=1339058 $Y=1343730
X2988 26 391 12258 14133 14053 25 14150 14213 14222 396 418 13518 14338 14346 3920 ICV_28 $T=1351020 1310770 0 0 $X=1351018 $Y=1310518
X2989 26 433 12050 14449 14454 25 14465 14472 14449 13687 438 13746 14454 14686 3920 ICV_28 $T=1371260 1244350 0 0 $X=1371258 $Y=1244098
X2990 26 437 12110 14389 14455 25 14150 14455 14481 396 420 13736 14562 14498 3920 ICV_28 $T=1371260 1296010 1 0 $X=1371258 $Y=1292070
X2991 26 447 12258 14589 14591 25 14599 451 14589 396 420 14391 14591 14424 3920 ICV_28 $T=1385060 1332910 0 0 $X=1385058 $Y=1332658
X2992 26 450 12051 14619 14626 25 14607 14636 14619 396 14673 14502 14626 14744 3920 ICV_28 $T=1387360 1296010 0 0 $X=1387358 $Y=1295758
X2993 26 14639 12754 14794 14797 25 14518 14768 14794 14831 14596 14663 14797 14876 3920 ICV_28 $T=1405760 1155790 0 0 $X=1405758 $Y=1155538
X2994 26 473 14913 14935 14860 25 14284 14962 14968 14831 488 13734 15030 15045 3920 ICV_28 $T=1422320 1126270 1 0 $X=1422318 $Y=1122330
X2995 26 14639 13329 14959 14898 25 14607 14898 14973 14810 469 14466 15040 14780 3920 ICV_28 $T=1423240 1273870 0 0 $X=1423238 $Y=1273618
X2996 26 489 12258 15093 15108 25 14599 15125 15093 483 478 15035 15108 15198 3920 ICV_28 $T=1439340 1340290 1 0 $X=1439338 $Y=1336350
X2997 26 15131 14966 15312 15368 25 15353 15413 15417 14831 488 13734 15453 15517 3920 ICV_28 $T=1468320 1126270 1 0 $X=1468318 $Y=1122330
X2998 26 475 13405 15448 15450 25 15135 15462 15448 15340 486 13745 15450 15553 3920 ICV_28 $T=1472460 1236970 0 0 $X=1472458 $Y=1236718
X2999 26 15075 15427 15463 15379 25 15135 15476 15463 15340 491 13948 15379 15568 3920 ICV_28 $T=1474760 1244350 0 0 $X=1474758 $Y=1244098
X3000 26 15253 15427 15513 15514 25 15353 15455 15513 15340 499 14838 15514 15654 3920 ICV_28 $T=1478900 1222210 0 0 $X=1478898 $Y=1221958
X3001 26 529 14937 15542 15506 25 15225 15506 15554 15340 499 14195 15662 15651 3920 ICV_28 $T=1482580 1303390 1 0 $X=1482578 $Y=1299450
X3002 26 15253 15224 15603 15605 25 15292 15617 15603 15340 512 14581 15605 15739 3920 ICV_28 $T=1489020 1281250 1 0 $X=1489018 $Y=1277310
X3003 26 518 14929 15618 15632 25 15225 15645 15656 534 519 14546 15619 15728 3920 ICV_28 $T=1491320 1325530 1 0 $X=1491318 $Y=1321590
X3004 26 15313 14992 15610 15640 25 15358 15640 15659 15687 15692 14839 15767 15683 3920 ICV_28 $T=1492240 1170550 1 0 $X=1492238 $Y=1166610
X3005 26 15313 14993 15636 15642 25 15353 15637 15636 15687 15321 14544 15642 15772 3920 ICV_28 $T=1492240 1200070 1 0 $X=1492238 $Y=1196130
X3006 26 15439 15427 15811 15842 25 15631 15848 15811 15340 515 14496 15842 15917 3920 ICV_28 $T=1509260 1229590 0 0 $X=1509258 $Y=1229338
X3007 26 521 16197 16075 16178 25 15631 16214 16250 16011 477 14580 16318 16099 3920 ICV_28 $T=1544680 1259110 1 0 $X=1544678 $Y=1255170
X3008 10870 10832 10908 8951 10811 10871 25 11021 26 MXI4X1 $T=1168400 1155790 1 0 $X=1168398 $Y=1151850
X3009 11102 10963 10908 8951 10756 10871 25 10867 26 MXI4X1 $T=1177140 1133650 0 180 $X=1168400 $Y=1129710
X3010 10878 10776 10908 8951 10772 10871 25 11173 26 MXI4X1 $T=1168860 1170550 0 0 $X=1168858 $Y=1170298
X3011 11031 10947 10908 8951 10901 10871 25 11201 26 MXI4X1 $T=1177140 1141030 0 0 $X=1177138 $Y=1140778
X3012 11054 10753 10908 8951 10984 10871 25 11226 26 MXI4X1 $T=1178060 1163170 1 0 $X=1178058 $Y=1159230
X3013 11107 10931 10908 8951 11067 10871 25 11261 26 MXI4X1 $T=1180360 1148410 0 0 $X=1180358 $Y=1148158
X3014 11303 10853 10908 11120 11125 141 25 11198 26 MXI4X1 $T=1193700 1177930 0 180 $X=1184960 $Y=1173990
X3015 11212 10946 10908 8951 11176 10871 25 11269 26 MXI4X1 $T=1185880 1126270 0 0 $X=1185878 $Y=1126018
X3016 11125 11120 10908 8951 10853 10871 25 11373 26 MXI4X1 $T=1185880 1170550 0 0 $X=1185878 $Y=1170298
X3017 13779 13807 352 13558 13804 359 25 13918 26 MXI4X1 $T=1316520 1296010 0 0 $X=1316518 $Y=1295758
X3018 13748 13761 354 13740 13824 13883 25 13920 26 MXI4X1 $T=1317900 1303390 0 0 $X=1317898 $Y=1303138
X3019 13779 13807 13853 13558 13804 364 25 14019 26 MXI4X1 $T=1320200 1296010 1 0 $X=1320198 $Y=1292070
X3020 13720 13754 13879 13769 13763 368 25 13926 26 MXI4X1 $T=1322960 1155790 1 0 $X=1322958 $Y=1151850
X3021 13859 13460 13880 13317 13755 369 25 13927 26 MXI4X1 $T=1322960 1163170 0 0 $X=1322958 $Y=1162918
X3022 13860 13877 13879 13557 13894 370 25 13928 26 MXI4X1 $T=1322960 1170550 1 0 $X=1322958 $Y=1166610
X3023 13868 13659 13879 13852 13907 364 25 13943 26 MXI4X1 $T=1323880 1133650 1 0 $X=1323878 $Y=1129710
X3024 13720 13754 13891 13769 13763 373 25 13966 26 MXI4X1 $T=1323880 1148410 0 0 $X=1323878 $Y=1148158
X3025 13869 13785 360 13561 13882 375 25 13949 26 MXI4X1 $T=1323880 1266490 0 0 $X=1323878 $Y=1266238
X3026 13869 13785 361 13561 13882 376 25 13957 26 MXI4X1 $T=1323880 1273870 1 0 $X=1323878 $Y=1269930
X3027 13844 13630 361 13655 13895 377 25 13972 26 MXI4X1 $T=1323880 1281250 1 0 $X=1323878 $Y=1277310
X3028 13870 13888 13893 13765 13788 370 25 13973 26 MXI4X1 $T=1323880 1325530 1 0 $X=1323878 $Y=1321590
X3029 13871 13889 13893 13368 13749 378 25 13953 26 MXI4X1 $T=1323880 1332910 1 0 $X=1323878 $Y=1328970
X3030 13819 13904 365 13784 13775 385 25 13975 26 MXI4X1 $T=1326180 1236970 1 0 $X=1326178 $Y=1233030
X3031 13790 13767 13880 13580 13780 13974 25 13986 26 MXI4X1 $T=1327560 1148410 1 0 $X=1327558 $Y=1144470
X3032 13905 13886 354 13455 13793 370 25 14018 26 MXI4X1 $T=1328020 1259110 1 0 $X=1328018 $Y=1255170
X3033 13819 13904 374 13784 13775 388 25 14017 26 MXI4X1 $T=1328940 1229590 0 0 $X=1328938 $Y=1229338
X3034 13905 13886 381 13455 13793 377 25 14033 26 MXI4X1 $T=1329860 1259110 0 0 $X=1329858 $Y=1258858
X3035 13748 13761 381 13740 13824 13974 25 14031 26 MXI4X1 $T=1329860 1310770 1 0 $X=1329858 $Y=1306830
X3036 13929 13637 360 13792 13963 368 25 14048 26 MXI4X1 $T=1331240 1251730 0 0 $X=1331238 $Y=1251478
X3037 13790 13767 13915 13580 13780 370 25 14055 26 MXI4X1 $T=1331700 1155790 1 0 $X=1331698 $Y=1151850
X3038 13753 13962 13880 14008 14001 389 25 14069 26 MXI4X1 $T=1333080 1141030 0 0 $X=1333078 $Y=1140778
X3039 13965 14009 365 13976 13945 385 25 14099 26 MXI4X1 $T=1334920 1236970 1 0 $X=1334918 $Y=1233030
X3040 13965 14009 374 13976 13945 373 25 14128 26 MXI4X1 $T=1338140 1229590 0 0 $X=1338138 $Y=1229338
X3041 13654 13954 13891 14039 13914 13974 25 14127 26 MXI4X1 $T=1338600 1126270 0 0 $X=1338598 $Y=1126018
X3042 14035 14058 360 14093 14103 398 25 14132 26 MXI4X1 $T=1338600 1259110 0 0 $X=1338598 $Y=1258858
X3043 13721 13592 13891 13723 13988 389 25 14171 26 MXI4X1 $T=1339060 1177930 0 0 $X=1339058 $Y=1177678
X3044 13654 13954 13879 14039 13914 364 25 14102 26 MXI4X1 $T=1339980 1133650 0 0 $X=1339978 $Y=1133398
X3045 14061 14060 354 14108 14114 13981 25 14138 26 MXI4X1 $T=1340440 1310770 1 0 $X=1340438 $Y=1306830
X3046 13721 13592 13879 13723 13988 398 25 14152 26 MXI4X1 $T=1340900 1185310 1 0 $X=1340898 $Y=1181370
X3047 13997 13916 14098 13816 14097 13974 25 14141 26 MXI4X1 $T=1340900 1214830 1 0 $X=1340898 $Y=1210890
X3048 13944 14101 13915 13995 14087 401 25 14151 26 MXI4X1 $T=1341820 1141030 0 0 $X=1341818 $Y=1140778
X3049 13944 14101 13880 13995 14087 376 25 14166 26 MXI4X1 $T=1342740 1141030 1 0 $X=1342738 $Y=1137090
X3050 13897 13341 14098 13791 14137 389 25 14205 26 MXI4X1 $T=1344120 1170550 1 0 $X=1344118 $Y=1166610
X3051 14126 14139 13912 14120 14182 389 25 14230 26 MXI4X1 $T=1346880 1332910 0 0 $X=1346878 $Y=1332658
X3052 14035 14058 361 14093 14103 369 25 14244 26 MXI4X1 $T=1347800 1259110 0 0 $X=1347798 $Y=1258858
X3053 14169 14172 361 14206 13923 415 25 14252 26 MXI4X1 $T=1351020 1281250 1 0 $X=1351018 $Y=1277310
X3054 14061 14060 381 14108 14114 388 25 14290 26 MXI4X1 $T=1351020 1310770 1 0 $X=1351018 $Y=1306830
X3055 13911 14154 13893 14153 14037 416 25 14259 26 MXI4X1 $T=1351020 1318150 0 0 $X=1351018 $Y=1317898
X3056 13911 14154 13912 14153 14037 415 25 14260 26 MXI4X1 $T=1351020 1325530 1 0 $X=1351018 $Y=1321590
X3057 14126 14139 13893 14120 14182 368 25 14261 26 MXI4X1 $T=1351020 1332910 1 0 $X=1351018 $Y=1328970
X3058 14168 14190 14119 14145 14220 368 25 14325 26 MXI4X1 $T=1352400 1207450 0 0 $X=1352398 $Y=1207198
X3059 14247 14256 13879 14186 14225 401 25 14143 26 MXI4X1 $T=1361140 1155790 0 180 $X=1352400 $Y=1151850
X3060 14168 14190 14098 14145 14220 359 25 14333 26 MXI4X1 $T=1352860 1214830 1 0 $X=1352858 $Y=1210890
X3061 13983 14210 365 14176 14187 13883 25 14242 26 MXI4X1 $T=1352860 1222210 0 0 $X=1352858 $Y=1221958
X3062 14173 14142 13853 14181 14212 416 25 14288 26 MXI4X1 $T=1352860 1288630 0 0 $X=1352858 $Y=1288378
X3063 14147 14146 14098 14091 14208 369 25 14351 26 MXI4X1 $T=1353780 1126270 0 0 $X=1353778 $Y=1126018
X3064 402 405 13853 403 419 416 25 14268 26 MXI4X1 $T=1354240 1347670 1 0 $X=1354238 $Y=1343730
X3065 14178 14184 371 14219 14298 389 25 14324 26 MXI4X1 $T=1357000 1192690 0 0 $X=1356998 $Y=1192438
X3066 14198 14250 354 14070 14216 398 25 14335 26 MXI4X1 $T=1357000 1251730 1 0 $X=1356998 $Y=1247790
X3067 14253 14235 13880 14214 14201 412 25 14231 26 MXI4X1 $T=1365740 1141030 0 180 $X=1357000 $Y=1137090
X3068 14178 14184 366 14219 14298 401 25 14353 26 MXI4X1 $T=1357920 1192690 1 0 $X=1357918 $Y=1188750
X3069 13983 14210 374 14176 14187 412 25 14292 26 MXI4X1 $T=1358380 1214830 0 0 $X=1358378 $Y=1214578
X3070 14255 14271 13879 14301 14315 368 25 14316 26 MXI4X1 $T=1358840 1148410 0 0 $X=1358838 $Y=1148158
X3071 14360 14337 360 14312 14299 14264 25 14227 26 MXI4X1 $T=1367580 1266490 0 180 $X=1358840 $Y=1262550
X3072 14198 14250 381 14070 14216 388 25 14385 26 MXI4X1 $T=1359300 1251730 0 0 $X=1359298 $Y=1251478
X3073 14255 14271 13891 14301 14315 376 25 14354 26 MXI4X1 $T=1359760 1148410 1 0 $X=1359758 $Y=1144470
X3074 14169 14172 360 14206 13923 385 25 14365 26 MXI4X1 $T=1359760 1281250 1 0 $X=1359758 $Y=1277310
X3075 13947 14096 14119 14285 14296 13883 25 14375 26 MXI4X1 $T=1360680 1163170 1 0 $X=1360678 $Y=1159230
X3076 14247 14256 13891 14186 14225 369 25 14237 26 MXI4X1 $T=1361140 1155790 1 0 $X=1361138 $Y=1151850
X3077 13947 14096 14098 14285 14296 386 25 14427 26 MXI4X1 $T=1364360 1170550 1 0 $X=1364358 $Y=1166610
X3078 14360 14337 361 14312 14299 13974 25 14317 26 MXI4X1 $T=1367580 1266490 1 0 $X=1367578 $Y=1262550
X3079 14484 14467 424 13984 14365 431 25 14240 26 MXI4X1 $T=1376780 1281250 1 180 $X=1368040 $Y=1280998
X3080 14491 14372 13893 14446 14424 13981 25 14341 26 MXI4X1 $T=1377700 1332910 1 180 $X=1368960 $Y=1332658
X3081 14493 14479 429 14116 14375 435 25 14380 26 MXI4X1 $T=1378160 1163170 0 180 $X=1369420 $Y=1159230
X3082 14494 14376 371 14453 14432 369 25 14257 26 MXI4X1 $T=1378160 1192690 0 180 $X=1369420 $Y=1188750
X3083 14436 14464 365 14239 14387 387 25 14144 26 MXI4X1 $T=1378620 1236970 0 180 $X=1369880 $Y=1233030
X3084 14498 14483 354 14438 14439 13883 25 14246 26 MXI4X1 $T=1378620 1288630 0 180 $X=1369880 $Y=1284690
X3085 14491 14372 13912 14446 14424 389 25 14319 26 MXI4X1 $T=1378620 1340290 0 180 $X=1369880 $Y=1336350
X3086 14475 14445 374 14418 14394 376 25 14355 26 MXI4X1 $T=1379080 1222210 1 180 $X=1370340 $Y=1221958
X3087 14498 14483 381 14438 14439 415 25 14358 26 MXI4X1 $T=1379080 1288630 1 180 $X=1370340 $Y=1288378
X3088 14540 14440 13880 14463 14433 389 25 14404 26 MXI4X1 $T=1380000 1141030 1 180 $X=1371260 $Y=1140778
X3089 14550 14510 13853 14346 14490 401 25 14357 26 MXI4X1 $T=1382760 1303390 0 180 $X=1374020 $Y=1299450
X3090 14540 14440 13915 14463 14433 416 25 14224 26 MXI4X1 $T=1383220 1148410 0 180 $X=1374480 $Y=1144470
X3091 14561 14524 361 14489 14501 13974 25 14318 26 MXI4X1 $T=1384140 1281250 0 180 $X=1375400 $Y=1277310
X3092 14550 14510 352 14346 14490 359 25 14331 26 MXI4X1 $T=1384140 1310770 0 180 $X=1375400 $Y=1306830
X3093 14553 14525 13893 14513 14503 368 25 14339 26 MXI4X1 $T=1384140 1318150 1 180 $X=1375400 $Y=1317898
X3094 14553 14525 13912 14513 14503 359 25 14340 26 MXI4X1 $T=1384140 1325530 0 180 $X=1375400 $Y=1321590
X3095 14547 14558 429 14179 14243 435 25 14495 26 MXI4X1 $T=1386900 1163170 0 180 $X=1378160 $Y=1159230
X3096 14494 14376 366 14453 14432 398 25 14474 26 MXI4X1 $T=1386900 1192690 0 180 $X=1378160 $Y=1188750
X3097 449 445 13853 443 442 375 25 14347 26 MXI4X1 $T=1386900 1347670 0 180 $X=1378160 $Y=1343730
X3098 14499 14556 371 14552 14539 369 25 14507 26 MXI4X1 $T=1387820 1207450 1 180 $X=1379080 $Y=1207198
X3099 14499 14556 366 14552 14539 364 25 14393 26 MXI4X1 $T=1384140 1200070 0 0 $X=1384138 $Y=1199818
X3100 14669 14638 14119 14611 14597 13883 25 14558 26 MXI4X1 $T=1393800 1155790 1 180 $X=1385060 $Y=1155538
X3101 14642 14571 14098 14595 14579 415 25 14555 26 MXI4X1 $T=1394260 1126270 1 180 $X=1385520 $Y=1126018
X3102 14669 14638 14098 14611 14597 13974 25 14523 26 MXI4X1 $T=1394260 1155790 0 180 $X=1385520 $Y=1151850
X3103 14567 14644 13915 14622 14604 13883 25 14479 26 MXI4X1 $T=1394260 1163170 1 180 $X=1385520 $Y=1162918
X3104 14707 14686 354 14677 14632 368 25 14476 26 MXI4X1 $T=1400240 1251730 0 180 $X=1391500 $Y=1247790
X3105 14736 14704 13893 14693 14678 370 25 14306 26 MXI4X1 $T=1401620 1318150 1 180 $X=1392880 $Y=1317898
X3106 14661 14590 14098 14628 14700 376 25 14664 26 MXI4X1 $T=1393800 1133650 1 0 $X=1393798 $Y=1129710
X3107 14688 14714 13891 14672 14687 13974 25 14215 26 MXI4X1 $T=1402540 1155790 1 180 $X=1393800 $Y=1155538
X3108 14715 14716 354 14699 14690 378 25 14437 26 MXI4X1 $T=1402540 1266490 1 180 $X=1393800 $Y=1266238
X3109 14661 14590 14119 14628 14700 13883 25 14493 26 MXI4X1 $T=1394260 1126270 0 0 $X=1394258 $Y=1126018
X3110 14688 14714 13879 14672 14687 458 25 14124 26 MXI4X1 $T=1403000 1155790 0 180 $X=1394260 $Y=1151850
X3111 14742 14710 14119 14702 14692 378 25 14367 26 MXI4X1 $T=1403000 1207450 1 180 $X=1394260 $Y=1207198
X3112 14742 14710 14098 14702 14692 388 25 14500 26 MXI4X1 $T=1407600 1214830 0 180 $X=1398860 $Y=1210890
X3113 14567 14644 13880 14622 14604 13974 25 14629 26 MXI4X1 $T=1399780 1170550 1 0 $X=1399778 $Y=1166610
X3114 14800 14783 13879 14774 14752 458 25 14291 26 MXI4X1 $T=1409440 1177930 1 180 $X=1400700 $Y=1177678
X3115 14740 14753 13853 14744 14784 375 25 14330 26 MXI4X1 $T=1402080 1296010 1 0 $X=1402078 $Y=1292070
X3116 14740 14753 352 14744 14784 359 25 14302 26 MXI4X1 $T=1402540 1296010 0 0 $X=1402538 $Y=1295758
X3117 14871 14813 360 14793 14780 387 25 14467 26 MXI4X1 $T=1412200 1273870 1 180 $X=1403460 $Y=1273618
X3118 14715 14716 381 14699 14690 377 25 14480 26 MXI4X1 $T=1404380 1273870 1 0 $X=1404378 $Y=1269930
X3119 14736 14704 13912 14693 14678 369 25 14307 26 MXI4X1 $T=1404380 1325530 1 0 $X=1404378 $Y=1321590
X3120 14800 14783 13891 14774 14752 388 25 14326 26 MXI4X1 $T=1413120 1177930 0 180 $X=1404380 $Y=1173990
X3121 14807 14788 371 14758 14757 13974 25 14286 26 MXI4X1 $T=1413120 1192690 1 180 $X=1404380 $Y=1192438
X3122 14812 14790 365 14745 14763 13883 25 14287 26 MXI4X1 $T=1413120 1229590 0 180 $X=1404380 $Y=1225650
X3123 14840 14818 381 14803 14789 369 25 14332 26 MXI4X1 $T=1413120 1303390 0 180 $X=1404380 $Y=1299450
X3124 14848 14689 374 14764 14791 412 25 14226 26 MXI4X1 $T=1413580 1236970 0 180 $X=1404840 $Y=1233030
X3125 14750 14776 13912 14785 14798 386 25 14295 26 MXI4X1 $T=1405760 1340290 0 0 $X=1405758 $Y=1340038
X3126 14876 14843 13880 14756 14811 412 25 14401 26 MXI4X1 $T=1415420 1141030 1 180 $X=1406680 $Y=1140778
X3127 14848 14689 365 14764 14791 14264 25 14125 26 MXI4X1 $T=1417260 1236970 1 180 $X=1408520 $Y=1236718
X3128 14876 14843 13915 14756 14811 364 25 14197 26 MXI4X1 $T=1418180 1141030 0 180 $X=1409440 $Y=1137090
X3129 468 471 13853 465 472 364 25 14313 26 MXI4X1 $T=1409900 1347670 0 0 $X=1409898 $Y=1347418
X3130 14884 14842 360 14857 14845 378 25 14199 26 MXI4X1 $T=1418640 1259110 0 180 $X=1409900 $Y=1255170
X3131 14884 14842 361 14857 14845 373 25 14293 26 MXI4X1 $T=1421860 1259110 1 180 $X=1413120 $Y=1258858
X3132 14787 14890 13880 14924 14893 386 25 14202 26 MXI4X1 $T=1418640 1148410 1 0 $X=1418638 $Y=1144470
X3133 14787 14890 13915 14924 14893 485 25 14107 26 MXI4X1 $T=1418640 1148410 0 0 $X=1418638 $Y=1148158
X3134 14975 14988 371 14995 14883 376 25 15065 26 MXI4X1 $T=1427840 1200070 0 0 $X=1427838 $Y=1199818
X3135 14975 14988 366 14995 14883 416 25 15059 26 MXI4X1 $T=1430140 1200070 1 0 $X=1430138 $Y=1196130
X3136 14978 15017 14098 15037 14974 369 25 15128 26 MXI4X1 $T=1432900 1170550 0 0 $X=1432898 $Y=1170298
X3137 15043 15025 381 15021 15048 388 25 15155 26 MXI4X1 $T=1437040 1266490 1 0 $X=1437038 $Y=1262550
X3138 15046 15063 14098 15039 15076 415 25 15143 26 MXI4X1 $T=1437500 1155790 1 0 $X=1437498 $Y=1151850
X3139 15046 15063 14119 15039 15076 385 25 15136 26 MXI4X1 $T=1437500 1155790 0 0 $X=1437498 $Y=1155538
X3140 14978 15017 14119 15037 14974 13883 25 15138 26 MXI4X1 $T=1437500 1170550 1 0 $X=1437498 $Y=1166610
X3141 15047 15018 366 14989 15077 13883 25 15140 26 MXI4X1 $T=1437500 1214830 0 0 $X=1437498 $Y=1214578
X3142 15043 15025 354 15021 15048 458 25 15141 26 MXI4X1 $T=1437500 1251730 0 0 $X=1437498 $Y=1251478
X3143 15049 15067 352 15072 14985 501 25 15142 26 MXI4X1 $T=1437500 1288630 0 0 $X=1437498 $Y=1288378
X3144 15049 15067 13853 15072 14985 364 25 15152 26 MXI4X1 $T=1438420 1288630 1 0 $X=1438418 $Y=1284690
X3145 15047 15018 371 14989 15077 501 25 15215 26 MXI4X1 $T=1438880 1214830 1 0 $X=1438878 $Y=1210890
X3146 15066 15082 371 15119 15127 388 25 15162 26 MXI4X1 $T=1439340 1200070 0 0 $X=1439338 $Y=1199818
X3147 15070 15088 13893 14940 15089 370 25 15220 26 MXI4X1 $T=1439800 1303390 0 0 $X=1439798 $Y=1303138
X3148 15190 15079 429 15136 15126 435 25 14543 26 MXI4X1 $T=1449000 1163170 1 180 $X=1440260 $Y=1162918
X3149 15070 15088 13912 14940 15089 388 25 15191 26 MXI4X1 $T=1440720 1310770 1 0 $X=1440718 $Y=1306830
X3150 15192 15160 14119 15139 15069 385 25 15079 26 MXI4X1 $T=1449920 1141030 0 180 $X=1441180 $Y=1137090
X3151 15106 15054 14119 15159 15045 13883 25 15204 26 MXI4X1 $T=1443940 1126270 1 0 $X=1443938 $Y=1122330
X3152 15106 15054 14098 15159 15045 415 25 15195 26 MXI4X1 $T=1444400 1126270 0 0 $X=1444398 $Y=1126018
X3153 15066 15082 366 15119 15127 416 25 15241 26 MXI4X1 $T=1444400 1200070 1 0 $X=1444398 $Y=1196130
X3154 15134 15151 13912 15166 15198 13974 25 15259 26 MXI4X1 $T=1444400 1332910 1 0 $X=1444398 $Y=1328970
X3155 498 502 13853 15061 15033 375 25 15230 26 MXI4X1 $T=1444400 1347670 1 0 $X=1444398 $Y=1343730
X3156 15228 15202 14119 15168 15161 385 25 15126 26 MXI4X1 $T=1453140 1163170 0 180 $X=1444400 $Y=1159230
X3157 15229 15204 429 15138 15148 435 25 14434 26 MXI4X1 $T=1453140 1170550 1 180 $X=1444400 $Y=1170298
X3158 15218 15150 381 15170 15163 373 25 15133 26 MXI4X1 $T=1453140 1251730 0 180 $X=1444400 $Y=1247790
X3159 15137 15157 13912 14934 15073 501 25 15227 26 MXI4X1 $T=1445320 1318150 0 0 $X=1445318 $Y=1317898
X3160 15228 15202 14098 15168 15161 412 25 15144 26 MXI4X1 $T=1454980 1155790 1 180 $X=1446240 $Y=1155538
X3161 15234 15216 14119 15203 15194 13883 25 15148 26 MXI4X1 $T=1454980 1170550 0 180 $X=1446240 $Y=1166610
X3162 498 502 352 15061 15033 501 25 508 26 MXI4X1 $T=1447620 1347670 0 0 $X=1447618 $Y=1347418
X3163 15221 15239 352 15265 15282 501 25 15297 26 MXI4X1 $T=1453140 1310770 1 0 $X=1453138 $Y=1306830
X3164 15221 15239 13853 15265 15282 485 25 15328 26 MXI4X1 $T=1453140 1310770 0 0 $X=1453138 $Y=1310518
X3165 15339 15281 13853 15219 15266 370 25 15208 26 MXI4X1 $T=1463720 1288630 0 180 $X=1454980 $Y=1284690
X3166 15339 15281 352 15219 15266 501 25 15233 26 MXI4X1 $T=1463720 1288630 1 180 $X=1454980 $Y=1288378
X3167 15234 15216 14098 15203 15194 13974 25 15217 26 MXI4X1 $T=1455900 1170550 1 0 $X=1455898 $Y=1166610
X3168 15360 15327 366 15322 15287 13883 25 15196 26 MXI4X1 $T=1464640 1214830 1 180 $X=1455900 $Y=1214578
X3169 15284 15288 366 15268 15252 13883 25 15149 26 MXI4X1 $T=1465100 1229590 0 180 $X=1456360 $Y=1225650
X3170 15330 15318 354 15280 15264 485 25 15231 26 MXI4X1 $T=1465100 1259110 0 180 $X=1456360 $Y=1255170
X3171 15192 15160 14098 15139 15069 373 25 15193 26 MXI4X1 $T=1459120 1141030 1 0 $X=1459118 $Y=1137090
X3172 15372 15354 352 15344 15319 501 25 509 26 MXI4X1 $T=1468320 1340290 1 180 $X=1459580 $Y=1340038
X3173 15325 15240 13880 15261 15356 373 25 15418 26 MXI4X1 $T=1461420 1148410 0 0 $X=1461418 $Y=1148158
X3174 15447 15375 366 15357 15317 375 25 15326 26 MXI4X1 $T=1470620 1200070 0 180 $X=1461880 $Y=1196130
X3175 15325 15240 13915 15261 15356 485 25 15419 26 MXI4X1 $T=1462800 1155790 0 0 $X=1462798 $Y=1155538
X3176 15411 15402 13853 15376 15363 416 25 15232 26 MXI4X1 $T=1472460 1288630 0 180 $X=1463720 $Y=1284690
X3177 15411 15402 352 15376 15363 501 25 15315 26 MXI4X1 $T=1472460 1288630 1 180 $X=1463720 $Y=1288378
X3178 15372 15354 13853 15344 15319 485 25 15333 26 MXI4X1 $T=1475220 1340290 0 180 $X=1466480 $Y=1336350
X3179 15447 15375 371 15357 15317 373 25 15256 26 MXI4X1 $T=1482120 1200070 1 180 $X=1473380 $Y=1199818
X3180 15484 15469 352 15442 15433 501 25 15336 26 MXI4X1 $T=1482120 1318150 1 180 $X=1473380 $Y=1317898
X3181 15432 15456 361 15361 15483 13974 25 15519 26 MXI4X1 $T=1473840 1281250 0 0 $X=1473838 $Y=1280998
X3182 15444 15466 360 15355 15488 14264 25 15522 26 MXI4X1 $T=1474760 1259110 0 0 $X=1474758 $Y=1258858
X3183 15432 15456 360 15361 15483 385 25 15544 26 MXI4X1 $T=1477980 1281250 1 0 $X=1477978 $Y=1277310
X3184 15480 15504 13879 15071 15531 13883 25 15563 26 MXI4X1 $T=1478900 1148410 0 0 $X=1478898 $Y=1148158
X3185 15482 15505 13915 15235 15528 398 25 15648 26 MXI4X1 $T=1478900 1185310 1 0 $X=1478898 $Y=1181370
X3186 15444 15466 361 15355 15488 386 25 15552 26 MXI4X1 $T=1478900 1266490 1 0 $X=1478898 $Y=1262550
X3187 15537 15407 13880 15409 15517 376 25 15478 26 MXI4X1 $T=1487640 1133650 0 180 $X=1478900 $Y=1129710
X3188 15558 15545 13891 15117 15521 373 25 15487 26 MXI4X1 $T=1488560 1192690 0 180 $X=1479820 $Y=1188750
X3189 15537 15407 13915 15409 15517 375 25 15510 26 MXI4X1 $T=1489940 1133650 1 180 $X=1481200 $Y=1133398
X3190 15480 15504 13891 15071 15531 389 25 15569 26 MXI4X1 $T=1482120 1148410 1 0 $X=1482118 $Y=1144470
X3191 15661 15643 424 15544 15606 52 25 14228 26 MXI4X1 $T=1497300 1281250 1 180 $X=1488560 $Y=1280998
X3192 15562 15464 13880 15612 15503 412 25 15641 26 MXI4X1 $T=1489020 1141030 1 0 $X=1489018 $Y=1137090
X3193 15555 15551 365 15526 15630 387 25 15665 26 MXI4X1 $T=1489020 1229590 0 0 $X=1489018 $Y=1229338
X3194 15377 15651 13912 15625 15609 412 25 15532 26 MXI4X1 $T=1497760 1310770 1 180 $X=1489020 $Y=1310518
X3195 15668 15652 13912 15626 15611 530 25 15534 26 MXI4X1 $T=1497760 1332910 0 180 $X=1489020 $Y=1328970
X3196 15558 15545 13879 15117 15521 458 25 15738 26 MXI4X1 $T=1489480 1185310 0 0 $X=1489478 $Y=1185058
X3197 15562 15464 13915 15612 15503 401 25 15672 26 MXI4X1 $T=1489940 1133650 0 0 $X=1489938 $Y=1133398
X3198 15668 15652 13893 15626 15611 13981 25 15539 26 MXI4X1 $T=1500060 1332910 1 180 $X=1491320 $Y=1332658
X3199 15555 15551 374 15526 15630 369 25 15752 26 MXI4X1 $T=1492240 1229590 1 0 $X=1492238 $Y=1225650
X3200 15628 15669 13891 15682 15713 13974 25 15721 26 MXI4X1 $T=1495920 1126270 0 0 $X=1495918 $Y=1126018
X3201 15628 15669 13879 15682 15713 13883 25 15679 26 MXI4X1 $T=1496380 1133650 1 0 $X=1496378 $Y=1129710
X3202 15629 15670 365 15688 15723 485 25 15735 26 MXI4X1 $T=1496380 1214830 0 0 $X=1496378 $Y=1214578
X3203 15751 15734 13879 15715 15683 13883 25 15658 26 MXI4X1 $T=1505120 1148410 1 180 $X=1496380 $Y=1148158
X3204 15803 15654 374 15716 15685 536 25 15653 26 MXI4X1 $T=1505120 1222210 1 180 $X=1496380 $Y=1221958
X3205 15754 15739 360 15724 15689 385 25 15643 26 MXI4X1 $T=1505580 1288630 0 180 $X=1496840 $Y=1284690
X3206 15754 15739 361 15724 15689 388 25 15667 26 MXI4X1 $T=1506040 1281250 1 180 $X=1497300 $Y=1280998
X3207 15766 15741 13912 15728 15695 537 25 15560 26 MXI4X1 $T=1506040 1340290 0 180 $X=1497300 $Y=1336350
X3208 15629 15670 374 15688 15723 412 25 15747 26 MXI4X1 $T=1497760 1214830 1 0 $X=1497758 $Y=1210890
X3209 15377 15651 13893 15625 15609 13981 25 15644 26 MXI4X1 $T=1497760 1310770 0 0 $X=1497758 $Y=1310518
X3210 15770 15635 13891 15729 15714 415 25 15655 26 MXI4X1 $T=1506500 1141030 0 180 $X=1497760 $Y=1137090
X3211 15756 15742 360 15732 15717 14264 25 15624 26 MXI4X1 $T=1506500 1266490 1 180 $X=1497760 $Y=1266238
X3212 15766 15741 13893 15728 15695 375 25 15573 26 MXI4X1 $T=1506500 1332910 0 180 $X=1497760 $Y=1328970
X3213 15773 15755 13893 15740 15727 416 25 15674 26 MXI4X1 $T=1507420 1303390 1 180 $X=1498680 $Y=1303138
X3214 15751 15734 13891 15715 15683 388 25 15677 26 MXI4X1 $T=1507880 1155790 1 180 $X=1499140 $Y=1155538
X3215 15568 15576 365 15553 15597 364 25 15761 26 MXI4X1 $T=1499600 1244350 1 0 $X=1499598 $Y=1240410
X3216 15753 15772 13891 15790 15805 412 25 15710 26 MXI4X1 $T=1505120 1192690 1 0 $X=1505118 $Y=1188750
X3217 15803 15654 365 15716 15685 13883 25 15748 26 MXI4X1 $T=1515240 1229590 0 180 $X=1506500 $Y=1225650
X3218 15753 15772 13879 15790 15805 370 25 15765 26 MXI4X1 $T=1507880 1185310 0 0 $X=1507878 $Y=1185058
X3219 15773 15755 13912 15740 15727 373 25 15559 26 MXI4X1 $T=1507880 1303390 0 0 $X=1507878 $Y=1303138
X3220 15850 15836 13915 15799 15784 375 25 15547 26 MXI4X1 $T=1516620 1155790 1 180 $X=1507880 $Y=1155538
X3221 15917 15880 553 15864 15858 14264 25 15780 26 MXI4X1 $T=1520760 1244350 0 180 $X=1512020 $Y=1240410
X3222 15775 15757 13880 15867 15879 412 25 15673 26 MXI4X1 $T=1513400 1170550 0 0 $X=1513398 $Y=1170298
X3223 15809 15860 361 15868 15881 376 25 15859 26 MXI4X1 $T=1513400 1273870 1 0 $X=1513398 $Y=1269930
X3224 15826 15887 374 15875 15863 386 25 15778 26 MXI4X1 $T=1522140 1222210 0 180 $X=1513400 $Y=1218270
X3225 15917 15880 554 15864 15858 376 25 15680 26 MXI4X1 $T=1522140 1236970 1 180 $X=1513400 $Y=1236718
X3226 15938 15869 554 15882 15861 550 25 15851 26 MXI4X1 $T=1522600 1288630 0 180 $X=1513860 $Y=1284690
X3227 15775 15757 13915 15867 15879 485 25 15771 26 MXI4X1 $T=1515240 1177930 0 0 $X=1515238 $Y=1177678
X3228 15826 15887 365 15875 15863 485 25 15789 26 MXI4X1 $T=1523980 1229590 0 180 $X=1515240 $Y=1225650
X3229 15809 15860 360 15868 15881 458 25 15664 26 MXI4X1 $T=1515700 1266490 0 0 $X=1515698 $Y=1266238
X3230 15938 15869 553 15882 15861 14264 25 15606 26 MXI4X1 $T=1525360 1281250 1 180 $X=1516620 $Y=1280998
X3231 118 25 9404 26 CLKINVX12 $T=1151840 1251730 1 0 $X=1151838 $Y=1247790
X3232 118 25 10868 26 CLKINVX12 $T=1211640 1296010 1 0 $X=1211638 $Y=1292070
X3233 12444 25 11826 26 CLKINVX12 $T=1245220 1177930 0 0 $X=1245218 $Y=1177678
X3234 13676 25 12746 26 CLKINVX12 $T=1304100 1303390 1 0 $X=1304098 $Y=1299450
X3235 12444 25 13599 26 CLKINVX12 $T=1348720 1133650 0 0 $X=1348718 $Y=1133398
X3236 13676 25 13687 26 CLKINVX12 $T=1358380 1244350 0 0 $X=1358378 $Y=1244098
X3237 12444 25 13998 26 CLKINVX12 $T=1374480 1170550 0 0 $X=1374478 $Y=1170298
X3238 13676 25 14810 26 CLKINVX12 $T=1449000 1288630 1 0 $X=1448998 $Y=1284690
X3239 15158 25 14865 26 CLKINVX12 $T=1450840 1207450 1 0 $X=1450838 $Y=1203510
X3240 15158 25 14831 26 CLKINVX12 $T=1453140 1141030 1 0 $X=1453138 $Y=1137090
X3241 15374 25 15340 26 CLKINVX12 $T=1495920 1266490 1 0 $X=1495918 $Y=1262550
X3242 15374 25 534 26 CLKINVX12 $T=1530420 1340290 1 0 $X=1530418 $Y=1336350
X3243 15158 25 15687 26 CLKINVX12 $T=1537780 1170550 1 0 $X=1537778 $Y=1166610
X3244 15374 25 16011 26 CLKINVX12 $T=1593900 1229590 0 0 $X=1593898 $Y=1229338
X3245 15374 25 595 26 CLKINVX12 $T=1597120 1340290 0 0 $X=1597118 $Y=1340038
X3246 14063 14055 59 14107 14123 399 26 25 14140 MX4X1 $T=1340900 1148410 0 0 $X=1340898 $Y=1148158
X3247 14102 13928 59 14124 14143 399 26 25 14174 MX4X1 $T=1343660 1155790 1 0 $X=1343658 $Y=1151850
X3248 14099 13975 59 14125 14144 399 26 25 14175 MX4X1 $T=1343660 1236970 1 0 $X=1343658 $Y=1233030
X3249 14151 13926 59 14197 14224 399 26 25 14248 MX4X1 $T=1350100 1148410 0 0 $X=1350098 $Y=1148158
X3250 14132 13949 59 14199 14227 52 26 25 14251 MX4X1 $T=1350100 1266490 1 0 $X=1350098 $Y=1262550
X3251 14069 13986 14191 14202 14231 78 26 25 14254 MX4X1 $T=1350560 1148410 1 0 $X=1350558 $Y=1144470
X3252 14127 13968 14191 14215 14237 410 26 25 14192 MX4X1 $T=1351940 1163170 1 0 $X=1351938 $Y=1159230
X3253 14128 14017 14191 14226 14245 410 26 25 14211 MX4X1 $T=1352400 1236970 1 0 $X=1352398 $Y=1233030
X3254 14138 13920 59 14229 14246 414 26 25 14272 MX4X1 $T=1352400 1303390 0 0 $X=1352398 $Y=1303138
X3255 14324 14011 422 14286 14257 413 26 25 14232 MX4X1 $T=1364820 1200070 0 180 $X=1356080 $Y=1196130
X3256 14242 14048 59 14287 14310 399 26 25 14329 MX4X1 $T=1357920 1229590 1 0 $X=1357918 $Y=1225650
X3257 13943 14152 59 14291 14316 399 26 25 14352 MX4X1 $T=1358380 1177930 0 0 $X=1358378 $Y=1177678
X3258 14244 13957 60 14293 14317 413 26 25 14305 MX4X1 $T=1358380 1266490 0 0 $X=1358378 $Y=1266238
X3259 14252 13972 60 14294 14318 413 26 25 14194 MX4X1 $T=1358380 1281250 0 0 $X=1358378 $Y=1280998
X3260 14230 14015 421 14295 14319 426 26 25 14371 MX4X1 $T=1358380 1332910 0 0 $X=1358378 $Y=1332658
X3261 14258 13918 421 14302 14331 426 26 25 14366 MX4X1 $T=1359300 1296010 0 0 $X=1359298 $Y=1295758
X3262 14259 13973 423 14306 14339 414 26 25 14359 MX4X1 $T=1359760 1318150 0 0 $X=1359758 $Y=1317898
X3263 14260 14000 421 14307 14340 426 26 25 14379 MX4X1 $T=1359760 1325530 1 0 $X=1359758 $Y=1321590
X3264 14261 13953 424 14309 14341 414 26 25 14361 MX4X1 $T=1359760 1332910 1 0 $X=1359758 $Y=1328970
X3265 14268 13991 59 14313 14347 414 26 25 14265 MX4X1 $T=1360220 1340290 0 0 $X=1360218 $Y=1340038
X3266 14025 14171 14191 14326 14354 413 26 25 14392 MX4X1 $T=1361600 1170550 0 0 $X=1361598 $Y=1170298
X3267 14292 14065 14191 14328 14355 78 26 25 14382 MX4X1 $T=1361600 1222210 0 0 $X=1361598 $Y=1221958
X3268 14288 14019 59 14330 14357 414 26 25 14388 MX4X1 $T=1361600 1288630 0 0 $X=1361598 $Y=1288378
X3269 14290 14031 421 14332 14358 426 26 25 14390 MX4X1 $T=1361600 1303390 1 0 $X=1361598 $Y=1299450
X3270 14325 14180 429 14367 14393 435 26 25 14441 MX4X1 $T=1364820 1207450 1 0 $X=1364818 $Y=1203510
X3271 14166 13966 14191 14401 14404 410 26 25 14478 MX4X1 $T=1367580 1148410 0 0 $X=1367578 $Y=1148158
X3272 14353 13989 429 14435 14474 435 26 25 14516 MX4X1 $T=1369880 1192690 0 0 $X=1369878 $Y=1192438
X3273 14335 14018 429 14437 14476 435 26 25 14517 MX4X1 $T=1369880 1251730 0 0 $X=1369878 $Y=1251478
X3274 14385 14033 422 14480 14497 78 26 25 14521 MX4X1 $T=1372640 1259110 0 0 $X=1372638 $Y=1258858
X3275 14333 14141 422 14500 14507 78 26 25 14570 MX4X1 $T=1375400 1214830 1 0 $X=1375398 $Y=1210890
X3276 14351 14205 422 14523 14555 426 26 25 14520 MX4X1 $T=1378620 1170550 1 0 $X=1378618 $Y=1166610
X3277 14427 13927 422 14629 14664 426 26 25 14566 MX4X1 $T=1387360 1170550 1 0 $X=1387358 $Y=1166610
X3278 15223 15155 422 15133 15121 78 26 25 14560 MX4X1 $T=1449000 1259110 0 180 $X=1440260 $Y=1255170
X3279 15196 15140 429 15149 15130 435 26 25 14386 MX4X1 $T=1449920 1222210 0 180 $X=1441180 $Y=1218270
X3280 15217 15128 422 15195 15156 413 26 25 14598 MX4X1 $T=1453140 1177930 0 180 $X=1444400 $Y=1173990
X3281 15144 15143 422 15193 15209 78 26 25 14559 MX4X1 $T=1446240 1155790 1 0 $X=1446238 $Y=1151850
X3282 15236 15215 422 15206 15169 78 26 25 14616 MX4X1 $T=1454980 1214830 1 180 $X=1446240 $Y=1214578
X3283 15231 15141 429 15207 15171 435 26 25 14554 MX4X1 $T=1454980 1251730 1 180 $X=1446240 $Y=1251478
X3284 15232 15152 59 15208 15172 414 26 25 14594 MX4X1 $T=1454980 1288630 1 180 $X=1446240 $Y=1288378
X3285 15256 15065 422 15162 15205 410 26 25 14322 MX4X1 $T=1456820 1200070 1 180 $X=1448080 $Y=1199818
X3286 15315 15142 421 15233 15211 426 26 25 14402 MX4X1 $T=1458200 1296010 0 180 $X=1449460 $Y=1292070
X3287 15326 15059 429 15241 15251 435 26 25 14565 MX4X1 $T=1461880 1192690 1 180 $X=1453140 $Y=1192438
X3288 15336 15227 421 15297 15269 426 26 25 14471 MX4X1 $T=1463260 1318150 1 180 $X=1454520 $Y=1317898
X3289 15347 15250 59 15328 15290 414 26 25 14383 MX4X1 $T=1465100 1325530 0 180 $X=1456360 $Y=1321590
X3290 507 15230 59 15333 15348 414 26 25 14241 MX4X1 $T=1459120 1347670 1 0 $X=1459118 $Y=1343730
X3291 15571 15418 14191 15478 15481 78 26 25 14369 MX4X1 $T=1484880 1155790 0 180 $X=1476140 $Y=1151850
X3292 15547 15419 59 15510 15511 399 26 25 14217 MX4X1 $T=1487180 1155790 1 180 $X=1478440 $Y=1155538
X3293 15559 15191 421 15532 15515 426 26 25 14450 MX4X1 $T=1487640 1310770 1 180 $X=1478900 $Y=1310518
X3294 15560 15259 421 15534 15516 426 26 25 14431 MX4X1 $T=1487640 1332910 0 180 $X=1478900 $Y=1328970
X3295 15573 15271 59 15539 15520 414 26 25 14308 MX4X1 $T=1488560 1332910 1 180 $X=1479820 $Y=1332658
X3296 15664 15522 424 15624 15598 52 26 25 14417 MX4X1 $T=1497300 1266490 1 180 $X=1488560 $Y=1266238
X3297 15673 15564 14191 15641 15614 78 26 25 14515 MX4X1 $T=1498680 1177930 0 180 $X=1489940 $Y=1173990
X3298 15674 15220 59 15644 15615 414 26 25 14350 MX4X1 $T=1498680 1303390 1 180 $X=1489940 $Y=1303138
X3299 15710 15487 14191 15655 15622 78 26 25 14218 MX4X1 $T=1499600 1192690 0 180 $X=1490860 $Y=1188750
X3300 15680 15666 14191 15653 15623 78 26 25 14236 MX4X1 $T=1499600 1236970 1 180 $X=1490860 $Y=1236718
X3301 15658 15563 59 15679 15660 399 26 25 14321 MX4X1 $T=1502820 1155790 0 180 $X=1494080 $Y=1151850
X3302 15677 15569 14191 15721 15678 78 26 25 14468 MX4X1 $T=1505120 1148410 0 180 $X=1496380 $Y=1144470
X3303 15765 15738 59 15675 15684 399 26 25 14207 MX4X1 $T=1505580 1185310 0 180 $X=1496840 $Y=1181370
X3304 15789 15665 59 15735 15693 399 26 25 14356 MX4X1 $T=1506500 1229590 1 180 $X=1497760 $Y=1229338
X3305 15771 15648 59 15672 15722 399 26 25 14342 MX4X1 $T=1507420 1177930 0 180 $X=1498680 $Y=1173990
X3306 15778 15752 14191 15747 15730 78 26 25 14430 MX4X1 $T=1508340 1222210 0 180 $X=1499600 $Y=1218270
X3307 15780 15761 59 15748 15731 399 26 25 14131 MX4X1 $T=1508340 1236970 1 180 $X=1499600 $Y=1236718
X3308 15851 15519 60 15667 15791 413 26 25 14221 MX4X1 $T=1514780 1281250 1 180 $X=1506040 $Y=1280998
X3309 15859 15552 60 15726 15800 413 26 25 14348 MX4X1 $T=1515700 1266490 1 180 $X=1506960 $Y=1266238
X3310 83 14254 11672 14369 25 26 MXI2X2 $T=1363900 1155790 0 0 $X=1363898 $Y=1155538
X3311 9371 35 26 25 INVX12 $T=1095720 1251730 1 180 $X=1092040 $Y=1251478
X3312 9721 65 26 25 INVX12 $T=1113200 1244350 0 180 $X=1109520 $Y=1240410
X3313 9763 73 26 25 INVX12 $T=1115040 1244350 1 180 $X=1111360 $Y=1244098
X3314 10063 97 26 25 INVX12 $T=1129760 1200070 1 180 $X=1126080 $Y=1199818
X3315 10075 94 26 25 INVX12 $T=1130220 1251730 0 180 $X=1126540 $Y=1247790
X3316 10039 101 26 25 INVX12 $T=1132060 1207450 0 0 $X=1132058 $Y=1207198
X3317 10238 108 26 25 INVX12 $T=1139420 1214830 0 0 $X=1139418 $Y=1214578
X3318 10350 113 26 25 INVX12 $T=1145860 1244350 1 0 $X=1145858 $Y=1240410
X3319 10580 119 26 25 INVX12 $T=1154140 1200070 1 0 $X=1154138 $Y=1196130
X3320 10715 123 26 25 INVX12 $T=1161500 1236970 0 180 $X=1157820 $Y=1233030
X3321 10765 127 26 25 INVX12 $T=1164720 1192690 0 180 $X=1161040 $Y=1188750
X3322 10767 133 26 25 INVX12 $T=1164720 1207450 0 180 $X=1161040 $Y=1203510
X3323 10768 128 26 25 INVX12 $T=1164720 1266490 1 180 $X=1161040 $Y=1266238
X3324 10734 130 26 25 INVX12 $T=1161500 1251730 1 0 $X=1161498 $Y=1247790
X3325 10789 132 26 25 INVX12 $T=1165640 1222210 0 180 $X=1161960 $Y=1218270
X3326 10790 135 26 25 INVX12 $T=1165640 1259110 1 180 $X=1161960 $Y=1258858
X3327 10808 131 26 25 INVX12 $T=1166560 1244350 0 180 $X=1162880 $Y=1240410
X3328 10829 136 26 25 INVX12 $T=1165640 1214830 0 0 $X=1165638 $Y=1214578
X3329 10960 145 26 25 INVX12 $T=1174840 1303390 1 180 $X=1171160 $Y=1303138
X3330 11104 154 26 25 INVX12 $T=1181280 1310770 0 180 $X=1177600 $Y=1306830
X3331 11123 155 26 25 INVX12 $T=1182200 1296010 0 180 $X=1178520 $Y=1292070
X3332 11059 157 26 25 INVX12 $T=1178980 1222210 1 0 $X=1178978 $Y=1218270
X3333 11129 152 26 25 INVX12 $T=1182660 1229590 1 180 $X=1178980 $Y=1229338
X3334 171 174 26 25 INVX12 $T=1188640 1288630 1 0 $X=1188638 $Y=1284690
X3335 11356 176 26 25 INVX12 $T=1192320 1310770 1 0 $X=1192318 $Y=1306830
X3336 11352 175 26 25 INVX12 $T=1206580 1207450 1 0 $X=1206578 $Y=1203510
X3337 316 323 26 25 INVX12 $T=1293060 1332910 1 0 $X=1293058 $Y=1328970
X3338 331 322 26 25 INVX12 $T=1299960 1244350 1 0 $X=1299958 $Y=1240410
X3339 510 258 26 25 INVX12 $T=1459580 1081990 1 0 $X=1459578 $Y=1078050
X3340 441 341 26 25 INVX12 $T=1476140 1104130 1 0 $X=1476138 $Y=1100190
X3341 457 540 26 25 INVX12 $T=1497300 1104130 0 0 $X=1497298 $Y=1103878
X3342 464 539 26 25 INVX12 $T=1499140 1089370 1 0 $X=1499138 $Y=1085430
X3343 14007 596 26 25 INVX12 $T=1564920 1163170 1 0 $X=1564918 $Y=1159230
X3344 615 617 26 25 INVX12 $T=1595740 1207450 1 0 $X=1595738 $Y=1203510
X3345 13684 645 26 25 INVX12 $T=1845520 1059850 0 0 $X=1845518 $Y=1059598
X3346 9428 9420 9481 26 25 9522 CLKMX2X2 $T=1097560 1229590 1 0 $X=1097558 $Y=1225650
X3347 9259 9525 9570 26 25 9593 CLKMX2X2 $T=1102160 1177930 0 0 $X=1102158 $Y=1177678
X3348 9680 9525 9570 26 25 9743 CLKMX2X2 $T=1109980 1177930 0 0 $X=1109978 $Y=1177678
X3349 9812 9525 9570 26 25 9600 CLKMX2X2 $T=1113660 1163170 1 180 $X=1109980 $Y=1162918
X3350 9775 57 64 26 25 9623 CLKMX2X2 $T=1114120 1318150 0 180 $X=1110440 $Y=1314210
X3351 9259 9713 9754 26 25 9885 CLKMX2X2 $T=1111360 1185310 1 0 $X=1111358 $Y=1181370
X3352 9884 9765 9667 26 25 9429 CLKMX2X2 $T=1115040 1126270 1 180 $X=1111360 $Y=1126018
X3353 9775 40 9660 26 25 9594 CLKMX2X2 $T=1115040 1251730 0 180 $X=1111360 $Y=1247790
X3354 9779 9729 9667 26 25 9685 CLKMX2X2 $T=1115500 1126270 0 180 $X=1111820 $Y=1122330
X3355 9836 9765 9667 26 25 9690 CLKMX2X2 $T=1118260 1148410 1 180 $X=1114580 $Y=1148158
X3356 9170 9525 9570 26 25 9895 CLKMX2X2 $T=1116880 1177930 0 0 $X=1116878 $Y=1177678
X3357 10057 9525 9570 26 25 9716 CLKMX2X2 $T=1123320 1148410 0 180 $X=1119640 $Y=1144470
X3358 9678 9525 9570 26 25 9790 CLKMX2X2 $T=1120560 1141030 1 0 $X=1120558 $Y=1137090
X3359 10061 9525 9570 26 25 9839 CLKMX2X2 $T=1124700 1163170 1 180 $X=1121020 $Y=1162918
X3360 10211 9525 9570 26 25 10072 CLKMX2X2 $T=1135280 1126270 0 180 $X=1131600 $Y=1122330
X3361 10185 10151 10221 26 25 10263 CLKMX2X2 $T=1133440 1096750 1 0 $X=1133438 $Y=1092810
X3362 10185 10221 10222 26 25 10288 CLKMX2X2 $T=1134820 1096750 0 0 $X=1134818 $Y=1096498
X3363 10185 10308 10246 26 25 10241 CLKMX2X2 $T=1140800 1074610 0 180 $X=1137120 $Y=1070670
X3364 10185 10309 10151 26 25 10257 CLKMX2X2 $T=1140800 1074610 1 180 $X=1137120 $Y=1074358
X3365 10332 9525 10216 26 25 10258 CLKMX2X2 $T=1140800 1148410 0 180 $X=1137120 $Y=1144470
X3366 10185 10246 10255 26 25 10398 CLKMX2X2 $T=1137580 1081990 1 0 $X=1137578 $Y=1078050
X3367 10266 10263 10192 26 25 10321 CLKMX2X2 $T=1137580 1104130 1 0 $X=1137578 $Y=1100190
X3368 10266 10241 10287 26 25 10124 CLKMX2X2 $T=1138040 1081990 0 0 $X=1138038 $Y=1081738
X3369 10412 9525 10216 26 25 10272 CLKMX2X2 $T=1141720 1155790 0 180 $X=1138040 $Y=1151850
X3370 10185 10414 10309 26 25 10464 CLKMX2X2 $T=1144020 1074610 0 0 $X=1144018 $Y=1074358
X3371 10266 10257 10288 26 25 10466 CLKMX2X2 $T=1144480 1111510 0 0 $X=1144478 $Y=1111258
X3372 10266 10463 10398 26 25 10393 CLKMX2X2 $T=1148160 1081990 0 180 $X=1144480 $Y=1078050
X3373 10185 10387 10308 26 25 10463 CLKMX2X2 $T=1145860 1067230 0 0 $X=1145858 $Y=1066978
X3374 10185 10489 10387 26 25 10432 CLKMX2X2 $T=1149540 1067230 0 180 $X=1145860 $Y=1063290
X3375 9952 9525 10216 26 25 10450 CLKMX2X2 $T=1153220 1163170 0 180 $X=1149540 $Y=1159230
X3376 10412 10520 10565 26 25 10625 CLKMX2X2 $T=1150000 1148410 0 0 $X=1149998 $Y=1148158
X3377 10185 10574 10414 26 25 10529 CLKMX2X2 $T=1153680 1074610 0 180 $X=1150000 $Y=1070670
X3378 10266 10576 10464 26 25 10490 CLKMX2X2 $T=1153680 1096750 0 180 $X=1150000 $Y=1092810
X3379 10266 10629 10432 26 25 10493 CLKMX2X2 $T=1157820 1081990 1 180 $X=1154140 $Y=1081738
X3380 10185 10603 10628 26 25 10629 CLKMX2X2 $T=1154600 1067230 0 0 $X=1154598 $Y=1066978
X3381 10185 10628 10489 26 25 10575 CLKMX2X2 $T=1158280 1067230 0 180 $X=1154600 $Y=1063290
X3382 9918 9525 10216 26 25 10637 CLKMX2X2 $T=1155520 1141030 0 0 $X=1155518 $Y=1140778
X3383 9952 10610 10647 26 25 10733 CLKMX2X2 $T=1155520 1163170 1 0 $X=1155518 $Y=1159230
X3384 10185 10671 10574 26 25 10576 CLKMX2X2 $T=1159660 1074610 1 180 $X=1155980 $Y=1074358
X3385 10266 10672 10575 26 25 10615 CLKMX2X2 $T=1159660 1081990 0 180 $X=1155980 $Y=1078050
X3386 9918 10746 10779 26 25 10822 CLKMX2X2 $T=1161960 1141030 1 0 $X=1161958 $Y=1137090
X3387 10185 10786 10603 26 25 10672 CLKMX2X2 $T=1166560 1067230 1 180 $X=1162880 $Y=1066978
X3388 10185 10793 10671 26 25 10656 CLKMX2X2 $T=1167020 1081990 0 180 $X=1163340 $Y=1078050
X3389 10185 10852 10745 26 25 10763 CLKMX2X2 $T=1168400 1096750 0 180 $X=1164720 $Y=1092810
X3390 10871 10776 10772 26 25 10803 CLKMX2X2 $T=1168860 1170550 1 180 $X=1165180 $Y=1170298
X3391 9775 10669 9493 26 25 11070 CLKMX2X2 $T=1171620 1244350 1 0 $X=1171618 $Y=1240410
X3392 10871 10753 10984 26 25 11262 CLKMX2X2 $T=1180360 1163170 0 0 $X=1180358 $Y=1162918
X3393 10871 10931 11067 26 25 11197 CLKMX2X2 $T=1180820 1148410 1 0 $X=1180818 $Y=1144470
X3394 10871 10946 11176 26 25 11196 CLKMX2X2 $T=1181740 1126270 0 0 $X=1181738 $Y=1126018
X3395 10907 10843 11214 26 25 11267 CLKMX2X2 $T=1183580 1273870 1 0 $X=1183578 $Y=1269930
X3396 169 10674 11296 26 25 11304 CLKMX2X2 $T=1188180 1318150 1 0 $X=1188178 $Y=1314210
X3397 10908 11207 11253 26 25 11321 CLKMX2X2 $T=1188640 1141030 1 0 $X=1188638 $Y=1137090
X3398 11382 11105 11379 26 25 11439 CLKMX2X2 $T=1195080 1059850 1 0 $X=1195078 $Y=1055910
X3399 10907 10648 11443 26 25 195 CLKMX2X2 $T=1196000 1214830 0 0 $X=1195998 $Y=1214578
X3400 10907 10769 11468 26 25 11492 CLKMX2X2 $T=1197840 1303390 0 0 $X=1197838 $Y=1303138
X3401 10907 10973 185 26 25 11579 CLKMX2X2 $T=1198300 1259110 1 0 $X=1198298 $Y=1255170
X3402 10907 10612 186 26 25 11333 CLKMX2X2 $T=1198300 1318150 1 0 $X=1198298 $Y=1314210
X3403 10907 11282 11516 26 25 11311 CLKMX2X2 $T=1199680 1273870 0 0 $X=1199678 $Y=1273618
X3404 184 11008 11528 26 25 11562 CLKMX2X2 $T=1200600 1229590 0 0 $X=1200598 $Y=1229338
X3405 10907 10849 11558 26 25 11575 CLKMX2X2 $T=1202440 1288630 0 0 $X=1202438 $Y=1288378
X3406 10907 10781 11581 26 25 11402 CLKMX2X2 $T=1203820 1251730 1 0 $X=1203818 $Y=1247790
X3407 11591 11621 11590 26 25 11446 CLKMX2X2 $T=1209340 1192690 0 180 $X=1205660 $Y=1188750
X3408 10907 10492 11622 26 25 188 CLKMX2X2 $T=1206120 1214830 1 0 $X=1206118 $Y=1210890
X3409 10907 10925 194 26 25 179 CLKMX2X2 $T=1206580 1325530 1 0 $X=1206578 $Y=1321590
X3410 11591 10807 10216 26 25 11660 CLKMX2X2 $T=1207040 1185310 1 0 $X=1207038 $Y=1181370
X3411 10907 10800 11646 26 25 11522 CLKMX2X2 $T=1207040 1229590 0 0 $X=1207038 $Y=1229338
X3412 10907 10956 11661 26 25 196 CLKMX2X2 $T=1207500 1288630 0 0 $X=1207498 $Y=1288378
X3413 191 10894 11672 26 25 11246 CLKMX2X2 $T=1207960 1244350 0 0 $X=1207958 $Y=1244098
X3414 10907 11009 11673 26 25 189 CLKMX2X2 $T=1207960 1259110 0 0 $X=1207958 $Y=1258858
X3415 10907 11415 11781 26 25 11819 CLKMX2X2 $T=1213020 1200070 1 0 $X=1213018 $Y=1196130
X3416 11382 11797 11566 26 25 11627 CLKMX2X2 $T=1216700 1089370 0 180 $X=1213020 $Y=1085430
X3417 10907 11430 11800 26 25 11504 CLKMX2X2 $T=1213480 1222210 1 0 $X=1213478 $Y=1218270
X3418 11828 10807 10216 26 25 11610 CLKMX2X2 $T=1217160 1177930 0 180 $X=1213480 $Y=1173990
X3419 11382 11629 11847 26 25 11656 CLKMX2X2 $T=1214860 1045090 0 0 $X=1214858 $Y=1044838
X3420 11382 11724 11794 26 25 11658 CLKMX2X2 $T=1218540 1067230 1 180 $X=1214860 $Y=1066978
X3421 11874 10807 10216 26 25 11917 CLKMX2X2 $T=1218080 1133650 1 0 $X=1218078 $Y=1129710
X3422 11828 11887 11914 26 25 11747 CLKMX2X2 $T=1218540 1170550 1 0 $X=1218538 $Y=1166610
X3423 11389 11656 11924 26 25 11565 CLKMX2X2 $T=1219000 1037710 1 0 $X=1218998 $Y=1033770
X3424 11389 11888 11464 26 25 11956 CLKMX2X2 $T=1219000 1081990 1 0 $X=1218998 $Y=1078050
X3425 11382 11933 11797 26 25 11888 CLKMX2X2 $T=1222680 1089370 0 180 $X=1219000 $Y=1085430
X3426 11874 12007 11968 26 25 11909 CLKMX2X2 $T=1226820 1141030 1 180 $X=1223140 $Y=1140778
X3427 11389 11657 12011 26 25 11607 CLKMX2X2 $T=1223600 1045090 0 0 $X=1223598 $Y=1044838
X3428 184 11442 12014 26 25 197 CLKMX2X2 $T=1223600 1192690 0 0 $X=1223598 $Y=1192438
X3429 11389 11537 11925 26 25 11912 CLKMX2X2 $T=1227280 1067230 1 180 $X=1223600 $Y=1066978
X3430 10907 10600 215 26 25 199 CLKMX2X2 $T=1224520 1340290 0 0 $X=1224518 $Y=1340038
X3431 11382 12053 11838 26 25 11958 CLKMX2X2 $T=1228200 1059850 1 180 $X=1224520 $Y=1059598
X3432 11382 12054 12003 26 25 11796 CLKMX2X2 $T=1228200 1074610 1 180 $X=1224520 $Y=1074358
X3433 11382 12012 11933 26 25 11739 CLKMX2X2 $T=1228200 1081990 1 180 $X=1224520 $Y=1081738
X3434 12013 10807 10216 26 25 11913 CLKMX2X2 $T=1228200 1155790 1 180 $X=1224520 $Y=1155538
X3435 11382 12003 12012 26 25 11925 CLKMX2X2 $T=1228660 1081990 0 180 $X=1224980 $Y=1078050
X3436 11382 12126 12113 26 25 11924 CLKMX2X2 $T=1233260 1045090 0 180 $X=1229580 $Y=1041150
X3437 184 11441 12146 26 25 216 CLKMX2X2 $T=1230040 1192690 1 0 $X=1230038 $Y=1188750
X3438 169 11312 223 26 25 12173 CLKMX2X2 $T=1230040 1347670 0 0 $X=1230038 $Y=1347418
X3439 10907 10557 12156 26 25 204 CLKMX2X2 $T=1230500 1325530 0 0 $X=1230498 $Y=1325278
X3440 10907 11840 12162 26 25 12062 CLKMX2X2 $T=1230960 1200070 0 0 $X=1230958 $Y=1199818
X3441 169 10641 12164 26 25 203 CLKMX2X2 $T=1230960 1303390 1 0 $X=1230958 $Y=1299450
X3442 169 11043 224 26 25 12256 CLKMX2X2 $T=1230960 1310770 1 0 $X=1230958 $Y=1306830
X3443 10907 10558 12165 26 25 210 CLKMX2X2 $T=1230960 1340290 1 0 $X=1230958 $Y=1336350
X3444 11382 11794 12054 26 25 11537 CLKMX2X2 $T=1234640 1067230 1 180 $X=1230960 $Y=1066978
X3445 12013 12136 12169 26 25 12261 CLKMX2X2 $T=1231420 1155790 0 0 $X=1231418 $Y=1155538
X3446 11382 11847 12126 26 25 11657 CLKMX2X2 $T=1235100 1045090 1 180 $X=1231420 $Y=1044838
X3447 12191 10807 10216 26 25 12066 CLKMX2X2 $T=1235100 1133650 0 180 $X=1231420 $Y=1129710
X3448 11382 12222 12174 26 25 12151 CLKMX2X2 $T=1236480 1059850 0 180 $X=1232800 $Y=1055910
X3449 11382 12174 12053 26 25 11940 CLKMX2X2 $T=1236480 1059850 1 180 $X=1232800 $Y=1059598
X3450 12214 10807 10216 26 25 12265 CLKMX2X2 $T=1235100 1148410 0 0 $X=1235098 $Y=1148158
X3451 184 12211 12255 26 25 12379 CLKMX2X2 $T=1235560 1192690 0 0 $X=1235558 $Y=1192438
X3452 169 11086 226 26 25 11993 CLKMX2X2 $T=1236020 1325530 0 0 $X=1236018 $Y=1325278
X3453 12285 10807 10216 26 25 12153 CLKMX2X2 $T=1240620 1133650 1 180 $X=1236940 $Y=1133398
X3454 11382 12113 12222 26 25 12011 CLKMX2X2 $T=1237400 1052470 1 0 $X=1237398 $Y=1048530
X3455 12285 12293 12334 26 25 12462 CLKMX2X2 $T=1239700 1141030 1 0 $X=1239698 $Y=1137090
X3456 12191 12304 12210 26 25 12461 CLKMX2X2 $T=1240160 1126270 0 0 $X=1240158 $Y=1126018
X3457 169 10456 12359 26 25 217 CLKMX2X2 $T=1241080 1296010 1 0 $X=1241078 $Y=1292070
X3458 184 11671 12368 26 25 11315 CLKMX2X2 $T=1241540 1200070 0 0 $X=1241538 $Y=1199818
X3459 229 11410 12369 26 25 12344 CLKMX2X2 $T=1241540 1229590 0 0 $X=1241538 $Y=1229338
X3460 184 10730 12392 26 25 12114 CLKMX2X2 $T=1242460 1236970 1 0 $X=1242458 $Y=1233030
X3461 169 11604 234 26 25 12297 CLKMX2X2 $T=1242920 1347670 1 0 $X=1242918 $Y=1343730
X3462 184 12118 12501 26 25 12303 CLKMX2X2 $T=1247060 1200070 1 0 $X=1247058 $Y=1196130
X3463 12214 12446 12438 26 25 12597 CLKMX2X2 $T=1247520 1148410 1 0 $X=1247518 $Y=1144470
X3464 229 12598 12651 26 25 236 CLKMX2X2 $T=1253500 1236970 1 0 $X=1253498 $Y=1233030
X3465 12678 12447 12719 26 25 12752 CLKMX2X2 $T=1256720 1148410 1 0 $X=1256718 $Y=1144470
X3466 229 12135 253 26 25 12803 CLKMX2X2 $T=1256720 1288630 1 0 $X=1256718 $Y=1284690
X3467 12863 10807 10216 26 25 12625 CLKMX2X2 $T=1261320 1170550 1 180 $X=1257640 $Y=1170298
X3468 184 12565 12758 26 25 12767 CLKMX2X2 $T=1258100 1192690 0 0 $X=1258098 $Y=1192438
X3469 12678 10807 10216 26 25 12709 CLKMX2X2 $T=1262240 1141030 1 180 $X=1258560 $Y=1140778
X3470 12815 10807 10216 26 25 12710 CLKMX2X2 $T=1262240 1163170 0 180 $X=1258560 $Y=1159230
X3471 169 12626 261 26 25 12835 CLKMX2X2 $T=1259940 1347670 1 0 $X=1259938 $Y=1343730
X3472 229 12652 12864 26 25 265 CLKMX2X2 $T=1263620 1273870 1 0 $X=1263618 $Y=1269930
X3473 12941 10807 10216 26 25 12854 CLKMX2X2 $T=1269140 1118890 1 180 $X=1265460 $Y=1118638
X3474 12863 12851 12920 26 25 12996 CLKMX2X2 $T=1265920 1177930 1 0 $X=1265918 $Y=1173990
X3475 229 12640 12921 26 25 246 CLKMX2X2 $T=1265920 1229590 1 0 $X=1265918 $Y=1225650
X3476 229 12195 12922 26 25 12694 CLKMX2X2 $T=1265920 1259110 0 0 $X=1265918 $Y=1258858
X3477 229 11484 271 26 25 13024 CLKMX2X2 $T=1265920 1303390 1 0 $X=1265918 $Y=1299450
X3478 229 12215 272 26 25 13025 CLKMX2X2 $T=1265920 1310770 1 0 $X=1265918 $Y=1306830
X3479 12955 10807 10216 26 25 12757 CLKMX2X2 $T=1269600 1126270 0 180 $X=1265920 $Y=1122330
X3480 12815 12931 12623 26 25 12862 CLKMX2X2 $T=1269600 1155790 1 180 $X=1265920 $Y=1155538
X3481 229 12503 274 26 25 12986 CLKMX2X2 $T=1266840 1281250 1 0 $X=1266838 $Y=1277310
X3482 229 12747 12946 26 25 244 CLKMX2X2 $T=1266840 1281250 0 0 $X=1266838 $Y=1280998
X3483 13010 10807 10216 26 25 12628 CLKMX2X2 $T=1270520 1126270 1 180 $X=1266840 $Y=1126018
X3484 12965 10807 10216 26 25 12882 CLKMX2X2 $T=1270520 1148410 0 180 $X=1266840 $Y=1144470
X3485 13065 10807 10216 26 25 12891 CLKMX2X2 $T=1270980 1170550 0 180 $X=1267300 $Y=1166610
X3486 13055 10807 10216 26 25 12942 CLKMX2X2 $T=1273740 1141030 0 180 $X=1270060 $Y=1137090
X3487 12955 13014 13059 26 25 13101 CLKMX2X2 $T=1271900 1118890 0 0 $X=1271898 $Y=1118638
X3488 13065 13113 12956 26 25 13023 CLKMX2X2 $T=1277880 1163170 1 180 $X=1274200 $Y=1162918
X3489 12965 13078 13112 26 25 13134 CLKMX2X2 $T=1274660 1148410 0 0 $X=1274658 $Y=1148158
X3490 229 12580 13114 26 25 13066 CLKMX2X2 $T=1274660 1236970 0 0 $X=1274658 $Y=1236718
X3491 13010 13015 13148 26 25 13111 CLKMX2X2 $T=1276040 1133650 1 0 $X=1276038 $Y=1129710
X3492 229 12335 13188 26 25 13183 CLKMX2X2 $T=1277420 1236970 1 0 $X=1277418 $Y=1233030
X3493 13055 13225 13241 26 25 13263 CLKMX2X2 $T=1281100 1141030 1 0 $X=1281098 $Y=1137090
X3494 229 12238 13300 26 25 12858 CLKMX2X2 $T=1283400 1259110 0 0 $X=1283398 $Y=1258858
X3495 12941 13303 13262 26 25 13123 CLKMX2X2 $T=1287080 1118890 1 180 $X=1283400 $Y=1118638
X3496 53 14240 14228 26 25 13300 CLKMX2X2 $T=1358380 1273870 1 180 $X=1354700 $Y=1273618
X3497 430 14380 14434 26 25 12162 CLKMX2X2 $T=1370800 1170550 0 0 $X=1370798 $Y=1170298
X3498 430 14495 14543 26 25 11781 CLKMX2X2 $T=1380920 1177930 1 0 $X=1380918 $Y=1173990
X3499 587 13628 16223 26 25 16339 CLKMX2X2 $T=1552960 1303390 1 0 $X=1552958 $Y=1299450
X3500 587 13811 16161 26 25 16329 CLKMX2X2 $T=1553420 1310770 0 0 $X=1553418 $Y=1310518
X3501 16519 16516 16435 26 25 14203 CLKMX2X2 $T=1575960 1266490 0 180 $X=1572280 $Y=1262550
X3502 603 601 16490 26 25 13471 CLKMX2X2 $T=1575960 1318150 0 180 $X=1572280 $Y=1314210
X3503 603 602 16491 26 25 13629 CLKMX2X2 $T=1575960 1347670 1 180 $X=1572280 $Y=1347418
X3504 603 605 16533 26 25 13811 CLKMX2X2 $T=1580100 1310770 1 180 $X=1576420 $Y=1310518
X3505 603 606 16526 26 25 13679 CLKMX2X2 $T=1580560 1347670 1 180 $X=1576880 $Y=1347418
X3506 603 16595 16534 26 25 276 CLKMX2X2 $T=1584240 1332910 0 180 $X=1580560 $Y=1328970
X3507 16519 609 16553 26 25 13628 CLKMX2X2 $T=1586540 1303390 0 180 $X=1582860 $Y=1299450
X3508 16519 16613 16583 26 25 13958 CLKMX2X2 $T=1588380 1229590 0 180 $X=1584700 $Y=1225650
X3509 16519 16628 16432 26 25 13567 CLKMX2X2 $T=1590680 1236970 1 180 $X=1587000 $Y=1236718
X3510 16519 611 16616 26 25 14743 CLKMX2X2 $T=1590680 1259110 0 180 $X=1587000 $Y=1255170
X3511 603 612 16617 26 25 13350 CLKMX2X2 $T=1590680 1318150 0 180 $X=1587000 $Y=1314210
X3512 16519 16634 16621 26 25 13843 CLKMX2X2 $T=1591140 1288630 0 180 $X=1587460 $Y=1284690
X3513 16519 16648 16566 26 25 13902 CLKMX2X2 $T=1592520 1229590 1 180 $X=1588840 $Y=1229338
X3514 16519 614 16629 26 25 13717 CLKMX2X2 $T=1592520 1303390 0 180 $X=1588840 $Y=1299450
X3515 16519 16650 16622 26 25 14833 CLKMX2X2 $T=1592980 1236970 0 180 $X=1589300 $Y=1233030
X3516 16519 16651 16623 26 25 13782 CLKMX2X2 $T=1592980 1244350 0 180 $X=1589300 $Y=1240410
X3517 16519 16652 16631 26 25 13881 CLKMX2X2 $T=1592980 1251730 0 180 $X=1589300 $Y=1247790
X3518 16519 16653 16633 26 25 13689 CLKMX2X2 $T=1592980 1266490 1 180 $X=1589300 $Y=1266238
X3519 16519 16654 16635 26 25 14741 CLKMX2X2 $T=1592980 1296010 1 180 $X=1589300 $Y=1295758
X3520 603 16712 16696 26 25 372 CLKMX2X2 $T=1598040 1318150 0 180 $X=1594360 $Y=1314210
X3521 603 16716 16675 26 25 325 CLKMX2X2 $T=1598500 1325530 1 180 $X=1594820 $Y=1325278
X3522 603 16725 16679 26 25 13235 CLKMX2X2 $T=1599880 1340290 0 180 $X=1596200 $Y=1336350
X3523 16519 16761 16698 26 25 13764 CLKMX2X2 $T=1602180 1229590 0 180 $X=1598500 $Y=1225650
X3524 603 626 16772 26 25 395 CLKMX2X2 $T=1608160 1340290 1 180 $X=1604480 $Y=1340038
X3525 603 16779 16773 26 25 330 CLKMX2X2 $T=1608620 1340290 0 180 $X=1604940 $Y=1336350
X3526 603 16782 16764 26 25 13786 CLKMX2X2 $T=1609540 1325530 1 180 $X=1605860 $Y=1325278
X3527 16519 16786 16780 26 25 14458 CLKMX2X2 $T=1610920 1251730 1 180 $X=1607240 $Y=1251478
X3528 16519 16787 16781 26 25 13725 CLKMX2X2 $T=1610920 1288630 0 180 $X=1607240 $Y=1284690
X3529 10207 25 26 10266 INVX2 $T=1153220 1089370 1 0 $X=1153218 $Y=1085430
X3530 11706 25 26 11744 INVX2 $T=1231420 1251730 1 0 $X=1231418 $Y=1247790
X3531 11736 25 26 11766 INVX2 $T=1232340 1259110 0 0 $X=1232338 $Y=1258858
X3532 14698 25 26 13942 INVX2 $T=1400700 1207450 1 0 $X=1400698 $Y=1203510
X3533 357 25 288 26 CLKINVX8 $T=1323880 1259110 0 0 $X=1323878 $Y=1258858
X3534 432 25 434 26 CLKINVX8 $T=1369420 1251730 1 0 $X=1369418 $Y=1247790
X3535 9283 26 8736 9300 25 NOR2XL $T=1088820 1192690 0 0 $X=1088818 $Y=1192438
X3536 9151 26 8948 9773 25 NOR2XL $T=1113200 1229590 1 0 $X=1113198 $Y=1225650
X3537 10002 26 9916 9734 25 NOR2XL $T=1122860 1111510 0 180 $X=1121480 $Y=1107570
X3538 9283 26 8881 10073 25 NOR2XL $T=1127460 1192690 0 0 $X=1127458 $Y=1192438
X3539 10136 26 9386 9858 25 NOR2XL $T=1133900 1081990 0 180 $X=1132520 $Y=1078050
X3540 10136 26 10435 10598 25 NOR2XL $T=1153220 1045090 0 0 $X=1153218 $Y=1044838
X3541 10404 26 134 10850 25 NOR2XL $T=1164720 1340290 0 0 $X=1164718 $Y=1340038
X3542 10770 26 134 137 25 NOR2XL $T=1165180 1347670 0 0 $X=1165178 $Y=1347418
X3543 10747 26 134 10876 25 NOR2XL $T=1166100 1340290 1 0 $X=1166098 $Y=1336350
X3544 10761 26 134 10961 25 NOR2XL $T=1168400 1332910 1 0 $X=1168398 $Y=1328970
X3545 10885 26 134 10880 25 NOR2XL $T=1170240 1340290 1 0 $X=1170238 $Y=1336350
X3546 10616 26 10445 11068 25 NOR2XL $T=1170700 1185310 0 0 $X=1170698 $Y=1185058
X3547 10889 26 134 10982 25 NOR2XL $T=1173920 1332910 0 0 $X=1173918 $Y=1332658
X3548 10380 26 11292 11332 25 NOR2XL $T=1190480 1259110 1 0 $X=1190478 $Y=1255170
X3549 10290 26 11336 11354 25 NOR2XL $T=1191860 1266490 1 0 $X=1191858 $Y=1262550
X3550 10122 26 11335 11306 25 NOR2XL $T=1193240 1185310 1 180 $X=1191860 $Y=1185058
X3551 11485 26 11242 11515 25 NOR2XL $T=1203820 1096750 1 180 $X=1202440 $Y=1096498
X3552 11587 26 11242 11717 25 NOR2XL $T=1207960 1096750 1 0 $X=1207958 $Y=1092810
X3553 11690 26 11242 11771 25 NOR2XL $T=1213940 1096750 1 0 $X=1213938 $Y=1092810
X3554 11383 26 11242 12292 25 NOR2XL $T=1231420 1089370 1 0 $X=1231418 $Y=1085430
X3555 12140 26 11242 12282 25 NOR2XL $T=1238320 1081990 1 0 $X=1238318 $Y=1078050
X3556 11846 26 11242 12254 25 NOR2XL $T=1238780 1045090 0 0 $X=1238778 $Y=1044838
X3557 12154 26 11023 12278 25 NOR2XL $T=1242460 1118890 0 180 $X=1241080 $Y=1114950
X3558 11763 26 11242 12690 25 NOR2XL $T=1242000 1037710 0 0 $X=1241998 $Y=1037458
X3559 11544 26 11242 12428 25 NOR2XL $T=1242460 1059850 1 0 $X=1242458 $Y=1055910
X3560 12048 26 11242 12443 25 NOR2XL $T=1242460 1059850 0 0 $X=1242458 $Y=1059598
X3561 11686 26 11242 12429 25 NOR2XL $T=1242460 1074610 1 0 $X=1242458 $Y=1070670
X3562 11218 26 11242 12450 25 NOR2XL $T=1242460 1074610 0 0 $X=1242458 $Y=1074358
X3563 11965 26 11242 12683 25 NOR2XL $T=1243380 1045090 0 0 $X=1243378 $Y=1044838
X3564 11294 26 11242 12402 25 NOR2XL $T=1243380 1067230 1 0 $X=1243378 $Y=1063290
X3565 12730 26 11225 12706 25 NOR2XL $T=1263160 1067230 1 180 $X=1261780 $Y=1066978
X3566 12880 26 12691 12829 25 NOR2XL $T=1267300 1089370 0 180 $X=1265920 $Y=1085430
X3567 12834 26 11295 13030 25 NOR2XL $T=1271900 1104130 0 0 $X=1271898 $Y=1103878
X3568 12154 26 11220 13554 25 NOR2XL $T=1296740 1141030 0 0 $X=1296738 $Y=1140778
X3569 8883 10055 26 25 10222 NOR2BXL $T=1132520 1104130 1 0 $X=1132518 $Y=1100190
X3570 11052 10470 26 25 11566 NOR2BXL $T=1203820 1089370 0 0 $X=1203818 $Y=1089118
X3571 12393 11323 26 25 12192 NOR2BXL $T=1245680 1170550 1 180 $X=1243840 $Y=1170298
X3572 9470 37 25 26 INVX3 $T=1096180 1310770 1 180 $X=1094800 $Y=1310518
X3573 9382 9504 25 26 INVX3 $T=1120100 1214830 1 0 $X=1120098 $Y=1210890
X3574 9382 9775 25 26 INVX3 $T=1123780 1214830 1 0 $X=1123778 $Y=1210890
X3575 10299 10185 25 26 INVX3 $T=1150460 1089370 1 0 $X=1150458 $Y=1085430
X3576 11030 11389 25 26 INVX3 $T=1196460 1037710 1 0 $X=1196458 $Y=1033770
X3577 11406 9196 25 26 INVX3 $T=1197840 1185310 0 180 $X=1196460 $Y=1181370
X3578 10951 11382 25 26 INVX3 $T=1209340 1045090 1 0 $X=1209338 $Y=1041150
X3579 492 25 12444 26 CLKBUFX16 $T=1438880 1236970 1 0 $X=1438878 $Y=1233030
X3580 8885 25 8748 8858 26 NAND2XL $T=1061680 1089370 1 180 $X=1060300 $Y=1089118
X3581 8917 25 8742 8939 26 NAND2XL $T=1063060 1074610 1 0 $X=1063058 $Y=1070670
X3582 9097 25 8871 9075 26 NAND2XL $T=1077320 1192690 0 180 $X=1075940 $Y=1188750
X3583 8885 25 8827 9110 26 NAND2XL $T=1076400 1074610 1 0 $X=1076398 $Y=1070670
X3584 9061 25 8749 9106 26 NAND2XL $T=1076400 1111510 0 0 $X=1076398 $Y=1111258
X3585 9110 25 9130 9115 26 NAND2XL $T=1077780 1067230 0 0 $X=1077778 $Y=1066978
X3586 9210 25 9227 9246 26 NAND2XL $T=1084680 1111510 1 0 $X=1084678 $Y=1107570
X3587 8834 25 8870 9241 26 NAND2XL $T=1086520 1074610 0 0 $X=1086518 $Y=1074358
X3588 8917 25 8822 9501 26 NAND2XL $T=1098480 1059850 0 0 $X=1098478 $Y=1059598
X3589 9283 25 8736 9332 26 NAND2XL $T=1100320 1192690 1 180 $X=1098940 $Y=1192438
X3590 9512 25 9228 9476 26 NAND2XL $T=1101700 1074610 1 0 $X=1101698 $Y=1070670
X3591 9238 25 9003 9339 26 NAND2XL $T=1104920 1111510 0 180 $X=1103540 $Y=1107570
X3592 9061 25 8880 9582 26 NAND2XL $T=1105840 1074610 1 0 $X=1105838 $Y=1070670
X3593 9138 25 9005 9621 26 NAND2XL $T=1105840 1074610 0 0 $X=1105838 $Y=1074358
X3594 8940 25 9624 9713 26 NAND2XL $T=1106300 1185310 0 0 $X=1106298 $Y=1185058
X3595 8948 25 9666 9619 26 NAND2XL $T=1110440 1229590 0 180 $X=1109060 $Y=1225650
X3596 8880 25 9708 9798 26 NAND2XL $T=1110900 1155790 1 0 $X=1110898 $Y=1151850
X3597 8870 25 9708 9859 26 NAND2XL $T=1111820 1170550 1 0 $X=1111818 $Y=1166610
X3598 9097 25 9006 9753 26 NAND2XL $T=1112280 1207450 1 0 $X=1112278 $Y=1203510
X3599 9258 25 9243 9835 26 NAND2XL $T=1115960 1067230 1 0 $X=1115958 $Y=1063290
X3600 9238 25 8980 9818 26 NAND2XL $T=1117800 1074610 0 0 $X=1117798 $Y=1074358
X3601 8822 25 9708 9989 26 NAND2XL $T=1121480 1141030 0 0 $X=1121478 $Y=1140778
X3602 8936 25 9708 10030 26 NAND2XL $T=1123320 1177930 0 0 $X=1123318 $Y=1177678
X3603 9509 25 9225 10080 26 NAND2XL $T=1128380 1185310 0 0 $X=1128378 $Y=1185058
X3604 8931 25 9708 10097 26 NAND2XL $T=1129300 1163170 0 0 $X=1129298 $Y=1162918
X3605 10080 25 10083 10138 26 NAND2XL $T=1129300 1185310 1 0 $X=1129298 $Y=1181370
X3606 10106 25 10124 10017 26 NAND2XL $T=1130220 1096750 1 0 $X=1130218 $Y=1092810
X3607 9283 25 8881 10109 26 NAND2XL $T=1132520 1192690 1 180 $X=1131140 $Y=1192438
X3608 10166 25 74 10032 26 NAND2XL $T=1133900 1303390 1 180 $X=1132520 $Y=1303138
X3609 9512 25 9437 10276 26 NAND2XL $T=1134820 1059850 1 0 $X=1134818 $Y=1055910
X3610 10106 25 10230 10120 26 NAND2XL $T=1135280 1111510 0 0 $X=1135278 $Y=1111258
X3611 10106 25 10321 10173 26 NAND2XL $T=1139880 1104130 0 0 $X=1139878 $Y=1103878
X3612 10353 25 104 10312 26 NAND2XL $T=1141720 1296010 1 180 $X=1140340 $Y=1295758
X3613 10106 25 10393 10037 26 NAND2XL $T=1145400 1104130 1 0 $X=1145398 $Y=1100190
X3614 10274 25 10337 10528 26 NAND2XL $T=1145400 1296010 1 0 $X=1145398 $Y=1292070
X3615 10472 25 10456 10307 26 NAND2XL $T=1147700 1281250 1 180 $X=1146320 $Y=1280998
X3616 10472 25 10557 10334 26 NAND2XL $T=1152760 1288630 0 180 $X=1151380 $Y=1284690
X3617 10472 25 10558 10148 26 NAND2XL $T=1152760 1296010 0 180 $X=1151380 $Y=1292070
X3618 10472 25 10600 10444 26 NAND2XL $T=1155520 1288630 1 180 $X=1154140 $Y=1288378
X3619 10472 25 10641 10572 26 NAND2XL $T=1158280 1296010 0 180 $X=1156900 $Y=1292070
X3620 10472 25 10648 10333 26 NAND2XL $T=1158740 1214830 1 180 $X=1157360 $Y=1214578
X3621 9806 25 10602 10564 26 NAND2XL $T=1158280 1052470 0 0 $X=1158278 $Y=1052218
X3622 10583 25 10732 10741 26 NAND2XL $T=1163800 1045090 0 180 $X=1162420 $Y=1041150
X3623 10472 25 10894 10611 26 NAND2XL $T=1170700 1236970 0 180 $X=1169320 $Y=1233030
X3624 10472 25 10925 10627 26 NAND2XL $T=1173000 1259110 0 180 $X=1171620 $Y=1255170
X3625 10472 25 10956 10146 26 NAND2XL $T=1174380 1281250 0 180 $X=1173000 $Y=1277310
X3626 10472 25 11008 10165 26 NAND2XL $T=1177140 1236970 1 180 $X=1175760 $Y=1236718
X3627 153 25 10982 11053 26 NAND2XL $T=1191400 1340290 0 180 $X=1190020 $Y=1336350
X3628 10972 25 11441 11121 26 NAND2XL $T=1199220 1200070 0 180 $X=1197840 $Y=1196130
X3629 10972 25 11442 10838 26 NAND2XL $T=1199220 1200070 1 180 $X=1197840 $Y=1199818
X3630 10972 25 11671 10839 26 NAND2XL $T=1212100 1200070 1 180 $X=1210720 $Y=1199818
X3631 11765 25 11740 11609 26 NAND2XL $T=1214860 1111510 1 180 $X=1213480 $Y=1111258
X3632 11839 25 11817 11687 26 NAND2XL $T=1217160 1118890 1 180 $X=1215780 $Y=1118638
X3633 11901 25 10967 11839 26 NAND2XL $T=1220380 1126270 1 180 $X=1219000 $Y=1126018
X3634 212 25 10876 11770 26 NAND2XL $T=1222220 1340290 1 180 $X=1220840 $Y=1340038
X3635 12236 25 12231 12149 26 NAND2XL $T=1236940 1118890 0 180 $X=1235560 $Y=1114950
X3636 12307 25 12267 12166 26 NAND2XL $T=1239700 1126270 0 180 $X=1238320 $Y=1122330
X3637 12363 25 12367 12145 26 NAND2XL $T=1244760 1111510 0 180 $X=1243380 $Y=1107570
X3638 12393 25 11323 12307 26 NAND2XL $T=1244760 1126270 0 180 $X=1243380 $Y=1122330
X3639 11926 25 11314 12391 26 NAND2XL $T=1243840 1163170 0 0 $X=1243838 $Y=1162918
X3640 12154 25 11023 12236 26 NAND2XL $T=1245680 1118890 0 180 $X=1244300 $Y=1114950
X3641 10972 25 237 12189 26 NAND2XL $T=1250280 1296010 0 180 $X=1248900 $Y=1292070
X3642 10972 25 239 12185 26 NAND2XL $T=1250740 1288630 1 180 $X=1249360 $Y=1288378
X3643 10972 25 240 11911 26 NAND2XL $T=1251660 1296010 1 180 $X=1250280 $Y=1295758
X3644 10972 25 12598 12675 26 NAND2XL $T=1252580 1229590 1 0 $X=1252578 $Y=1225650
X3645 10972 25 12640 12579 26 NAND2XL $T=1256260 1222210 1 180 $X=1254880 $Y=1221958
X3646 12714 25 12722 12180 26 NAND2XL $T=1260400 1052470 0 180 $X=1259020 $Y=1048530
X3647 10972 25 12747 12745 26 NAND2XL $T=1259480 1251730 1 0 $X=1259478 $Y=1247790
X3648 12500 25 11275 12363 26 NAND2XL $T=1260860 1111510 0 180 $X=1259480 $Y=1107570
X3649 10972 25 12652 12765 26 NAND2XL $T=1260400 1266490 1 0 $X=1260398 $Y=1262550
X3650 10972 25 259 12661 26 NAND2XL $T=1261780 1296010 0 180 $X=1260400 $Y=1292070
X3651 12685 25 11066 12714 26 NAND2XL $T=1262700 1059850 0 180 $X=1261320 $Y=1055910
X3652 10972 25 266 12816 26 NAND2XL $T=1266380 1244350 1 180 $X=1265000 $Y=1244098
X3653 12582 25 11063 12545 26 NAND2XL $T=1267300 1059850 0 180 $X=1265920 $Y=1055910
X3654 12750 25 12869 12715 26 NAND2XL $T=1267300 1067230 1 180 $X=1265920 $Y=1066978
X3655 12982 25 12870 12663 26 NAND2XL $T=1267300 1096750 0 180 $X=1265920 $Y=1092810
X3656 10972 25 269 12777 26 NAND2XL $T=1268680 1251730 0 180 $X=1267300 $Y=1247790
X3657 12744 25 9708 13014 26 NAND2XL $T=1267760 1118890 1 0 $X=1267758 $Y=1114950
X3658 12685 25 12889 12868 26 NAND2XL $T=1271900 1067230 1 0 $X=1271898 $Y=1063290
X3659 13104 25 13047 13035 26 NAND2XL $T=1274660 1052470 0 180 $X=1273280 $Y=1048530
X3660 12857 25 11087 12750 26 NAND2XL $T=1278340 1074610 1 180 $X=1276960 $Y=1074358
X3661 12943 25 11243 12982 26 NAND2XL $T=1279260 1089370 1 180 $X=1277880 $Y=1089118
X3662 13100 25 13147 12743 26 NAND2XL $T=1279260 1104130 1 180 $X=1277880 $Y=1103878
X3663 12929 25 11421 13100 26 NAND2XL $T=1280180 1111510 0 180 $X=1278800 $Y=1107570
X3664 12834 25 11295 12881 26 NAND2XL $T=1283860 1104130 1 180 $X=1282480 $Y=1103878
X3665 12926 25 9708 13303 26 NAND2XL $T=1282940 1118890 1 0 $X=1282938 $Y=1114950
X3666 12814 25 12874 13361 26 NAND2XL $T=1283400 1096750 0 0 $X=1283398 $Y=1096498
X3667 12857 25 12744 13232 26 NAND2XL $T=1285240 1074610 1 180 $X=1283860 $Y=1074358
X3668 12943 25 12927 13240 26 NAND2XL $T=1285240 1104130 1 0 $X=1285238 $Y=1100190
X3669 12393 25 11177 13427 26 NAND2XL $T=1289840 1141030 1 0 $X=1289838 $Y=1137090
X3670 12500 25 12463 13488 26 NAND2XL $T=1291220 1118890 0 0 $X=1291218 $Y=1118638
X3671 12929 25 13453 13459 26 NAND2XL $T=1293520 1104130 0 0 $X=1293518 $Y=1103878
X3672 13261 25 13463 13468 26 NAND2XL $T=1297200 1074610 1 180 $X=1295820 $Y=1074358
X3673 13546 25 13393 13446 26 NAND2XL $T=1297660 1089370 0 180 $X=1296280 $Y=1085430
X3674 13562 25 13586 13500 26 NAND2XL $T=1301340 1133650 0 180 $X=1299960 $Y=1129710
X3675 13474 25 13705 13709 26 NAND2XL $T=1310080 1111510 0 0 $X=1310078 $Y=1111258
X3676 8872 8947 25 8884 8951 26 9000 8999 OAI221XL $T=1067660 1170550 1 0 $X=1067658 $Y=1166610
X3677 8946 8827 25 8822 8872 26 9001 9011 OAI221XL $T=1067660 1170550 0 0 $X=1067658 $Y=1170298
X3678 9128 9086 25 9358 9242 26 9387 9402 OAI221XL $T=1093420 1133650 1 0 $X=1093418 $Y=1129710
X3679 9128 8966 25 9358 9467 26 9478 9684 OAI221XL $T=1097560 1126270 1 0 $X=1097558 $Y=1122330
X3680 8822 9353 25 9119 8936 26 9468 9658 OAI221XL $T=1103080 1141030 1 0 $X=1103078 $Y=1137090
X3681 10004 9922 25 9913 9897 26 9837 9848 OAI221XL $T=1123320 1273870 0 180 $X=1120100 $Y=1269930
X3682 10004 9994 25 9928 9897 26 9745 9524 OAI221XL $T=1124700 1281250 1 180 $X=1121480 $Y=1280998
X3683 10004 10050 25 9965 9897 26 9902 9616 OAI221XL $T=1125160 1251730 1 180 $X=1121940 $Y=1251478
X3684 10191 10095 25 10053 9897 26 9908 9975 OAI221XL $T=1129760 1236970 0 180 $X=1126540 $Y=1233030
X3685 10191 10074 25 10121 9897 26 10049 9993 OAI221XL $T=1132060 1244350 0 180 $X=1128840 $Y=1240410
X3686 10004 10248 25 10102 9897 26 10076 9617 OAI221XL $T=1132060 1273870 0 180 $X=1128840 $Y=1269930
X3687 10004 10265 25 10279 9897 26 9717 9523 OAI221XL $T=1139880 1259110 1 180 $X=1136660 $Y=1258858
X3688 10260 10121 25 10074 10290 26 10040 10310 OAI221XL $T=1137120 1244350 1 0 $X=1137118 $Y=1240410
X3689 10191 10296 25 10289 9897 26 10270 10237 OAI221XL $T=1140800 1207450 1 180 $X=1137580 $Y=1207198
X3690 10380 9913 25 9922 10290 26 10280 10231 OAI221XL $T=1141260 1266490 1 180 $X=1138040 $Y=1266238
X3691 10380 9965 25 10050 10290 26 10239 10297 OAI221XL $T=1142180 1259110 0 180 $X=1138960 $Y=1255170
X3692 10260 9928 25 9994 10281 26 10396 10413 OAI221XL $T=1141260 1288630 1 0 $X=1141258 $Y=1284690
X3693 10191 10571 25 10427 9897 26 10403 10031 OAI221XL $T=1146780 1222210 0 180 $X=1143560 $Y=1218270
X3694 10260 10102 25 10248 10290 26 10077 10409 OAI221XL $T=1147240 1273870 0 180 $X=1144020 $Y=1269930
X3695 10380 10480 25 10402 10426 26 10419 10382 OAI221XL $T=1147700 1207450 0 180 $X=1144480 $Y=1203510
X3696 10191 10454 25 10436 9897 26 10421 10156 OAI221XL $T=1147700 1244350 1 180 $X=1144480 $Y=1244098
X3697 10191 10402 25 10480 10373 26 10442 10361 OAI221XL $T=1149080 1200070 1 180 $X=1145860 $Y=1199818
X3698 10260 10053 25 10095 10290 26 10326 10364 OAI221XL $T=1149540 1229590 1 180 $X=1146320 $Y=1229338
X3699 10004 10546 25 10555 9897 26 10535 9361 OAI221XL $T=1153220 1273870 1 180 $X=1150000 $Y=1273618
X3700 10380 10289 25 10296 10426 26 10570 10556 OAI221XL $T=1150460 1207450 1 0 $X=1150458 $Y=1203510
X3701 10191 10588 25 10566 9897 26 10540 10351 OAI221XL $T=1153680 1251730 1 180 $X=1150460 $Y=1251478
X3702 10191 10626 25 10620 10373 26 10601 10401 OAI221XL $T=1157820 1200070 1 180 $X=1154600 $Y=1199818
X3703 10260 10279 25 10265 10290 26 10541 10640 OAI221XL $T=1155060 1259110 0 0 $X=1155058 $Y=1258858
X3704 10380 10620 25 10626 10426 26 10654 10673 OAI221XL $T=1155980 1207450 1 0 $X=1155978 $Y=1203510
X3705 10260 10555 25 10546 10290 26 10621 10617 OAI221XL $T=1159200 1273870 1 180 $X=1155980 $Y=1273618
X3706 10380 10436 25 10454 10290 26 10749 10758 OAI221XL $T=1160580 1244350 0 0 $X=1160578 $Y=1244098
X3707 10792 10004 25 10373 10743 26 10735 10543 OAI221XL $T=1164720 1303390 0 180 $X=1161500 $Y=1299450
X3708 10004 10791 25 10809 10373 26 10830 10841 OAI221XL $T=1164260 1296010 0 0 $X=1164258 $Y=1295758
X3709 10888 10004 25 10373 10840 26 10618 9738 OAI221XL $T=1169320 1288630 0 180 $X=1166100 $Y=1284690
X3710 10380 10427 25 10571 10426 26 10639 10893 OAI221XL $T=1167020 1222210 0 0 $X=1167018 $Y=1221958
X3711 10380 10566 25 10588 10290 26 10721 10813 OAI221XL $T=1170700 1251730 0 180 $X=1167480 $Y=1247790
X3712 10191 10919 25 10933 10373 26 10949 10959 OAI221XL $T=1171160 1229590 0 0 $X=1171158 $Y=1229338
X3713 10191 10766 25 10932 10373 26 10937 10996 OAI221XL $T=1172080 1200070 1 0 $X=1172078 $Y=1196130
X3714 10380 10932 25 10766 10426 26 10964 10953 OAI221XL $T=1172080 1200070 0 0 $X=1172078 $Y=1199818
X3715 9924 10445 25 10669 10147 26 10974 10988 OAI221XL $T=1172540 1273870 0 0 $X=1172538 $Y=1273618
X3716 10191 11114 25 11103 10373 26 10968 10950 OAI221XL $T=1181740 1266490 1 180 $X=1178520 $Y=1266238
X3717 10292 11111 25 11122 10373 26 11148 11252 OAI221XL $T=1180360 1288630 0 0 $X=1180358 $Y=1288378
X3718 10191 11085 25 11136 10373 26 11095 10997 OAI221XL $T=1183580 1200070 1 180 $X=1180360 $Y=1199818
X3719 10191 11202 25 11163 10373 26 11110 11041 OAI221XL $T=1184960 1259110 1 180 $X=1181740 $Y=1258858
X3720 10191 11266 25 11187 10373 26 11161 11154 OAI221XL $T=1186340 1207450 0 180 $X=1183120 $Y=1203510
X3721 10004 11216 25 11210 10373 26 11115 11024 OAI221XL $T=1187260 1303390 0 180 $X=1184040 $Y=1299450
X3722 10191 11230 25 11222 10373 26 11209 11022 OAI221XL $T=1188640 1229590 1 180 $X=1185420 $Y=1229338
X3723 10191 11336 25 11292 10373 26 11130 10905 OAI221XL $T=1191860 1251730 1 180 $X=1188640 $Y=1251478
X3724 10191 11310 25 11289 10373 26 11263 10981 OAI221XL $T=1192320 1214830 1 180 $X=1189100 $Y=1214578
X3725 10191 11374 25 11318 10373 26 11113 11006 OAI221XL $T=1193240 1244350 1 180 $X=1190020 $Y=1244098
X3726 10191 11285 25 11291 10373 26 11307 10941 OAI221XL $T=1194160 1236970 1 180 $X=1190940 $Y=1236718
X3727 10380 11136 25 11085 10426 26 11069 11357 OAI221XL $T=1197840 1200070 1 180 $X=1194620 $Y=1199818
X3728 10191 11465 25 11427 10373 26 11381 11239 OAI221XL $T=1199220 1222210 1 180 $X=1196000 $Y=1221958
X3729 10004 11431 25 11419 10373 26 11277 11240 OAI221XL $T=1200140 1303390 0 180 $X=1196920 $Y=1299450
X3730 10380 11427 25 11465 10426 26 11204 11728 OAI221XL $T=1201980 1222210 1 0 $X=1201978 $Y=1218270
X3731 11568 11451 25 11586 11563 26 11615 11624 OAI221XL $T=1205660 1310770 1 0 $X=1205658 $Y=1306830
X3732 11568 11542 25 11586 10220 26 11655 11769 OAI221XL $T=1207500 1303390 1 0 $X=1207498 $Y=1299450
X3733 11568 11633 25 11586 10942 26 11689 11623 OAI221XL $T=1208420 1266490 1 0 $X=1208418 $Y=1262550
X3734 11568 11625 25 11586 9803 26 11735 11793 OAI221XL $T=1211180 1310770 0 0 $X=1211178 $Y=1310518
X3735 11568 11688 25 11586 10999 26 11745 11843 OAI221XL $T=1211640 1251730 1 0 $X=1211638 $Y=1247790
X3736 11568 11645 25 11586 9827 26 11746 11757 OAI221XL $T=1211640 1273870 0 0 $X=1211638 $Y=1273618
X3737 11706 11729 25 11736 9827 26 11768 11784 OAI221XL $T=1212560 1281250 1 0 $X=1212558 $Y=1277310
X3738 11568 11705 25 11586 10485 26 11812 11758 OAI221XL $T=1213940 1288630 1 0 $X=1213938 $Y=1284690
X3739 11626 11752 25 11731 9803 26 11814 11830 OAI221XL $T=1213940 1318150 0 0 $X=1213938 $Y=1317898
X3740 11568 11674 25 11586 11827 26 11842 11904 OAI221XL $T=1214860 1236970 0 0 $X=1214858 $Y=1236718
X3741 11706 11756 25 11736 10999 26 11844 11872 OAI221XL $T=1214860 1251730 0 0 $X=1214858 $Y=1251478
X3742 11706 11779 25 11736 11071 26 11845 11873 OAI221XL $T=1214860 1266490 1 0 $X=1214858 $Y=1262550
X3743 11706 11967 25 11736 10485 26 11813 11787 OAI221XL $T=1219000 1288630 1 180 $X=1215780 $Y=1288378
X3744 11568 11734 25 11586 11071 26 11910 11906 OAI221XL $T=1218540 1259110 1 0 $X=1218538 $Y=1255170
X3745 11568 11903 25 11586 11810 26 11938 11971 OAI221XL $T=1219920 1207450 1 0 $X=1219918 $Y=1203510
X3746 11568 11918 25 11586 11896 26 11999 11981 OAI221XL $T=1223140 1214830 0 0 $X=1223138 $Y=1214578
X3747 11568 12106 25 11586 11932 26 11966 11959 OAI221XL $T=1226360 1236970 0 180 $X=1223140 $Y=1233030
X3748 11706 12010 25 11736 10220 26 11972 11864 OAI221XL $T=1226820 1303390 0 180 $X=1223600 $Y=1299450
X3749 11706 12137 25 11736 10942 26 12115 11767 OAI221XL $T=1233720 1273870 0 180 $X=1230500 $Y=1269930
X3750 11706 225 25 11736 11635 26 12239 12246 OAI221XL $T=1234180 1310770 0 0 $X=1234178 $Y=1310518
X3751 11706 12139 25 11736 12193 26 12257 12294 OAI221XL $T=1236020 1222210 0 0 $X=1236018 $Y=1221958
X3752 12270 12240 25 12296 11635 26 12271 12470 OAI221XL $T=1238780 1318150 1 0 $X=1238778 $Y=1314210
X3753 12270 12315 25 12296 12186 26 12348 12346 OAI221XL $T=1240620 1244350 0 0 $X=1240618 $Y=1244098
X3754 11568 12404 25 12296 12163 26 12331 12324 OAI221XL $T=1244760 1207450 1 180 $X=1241540 $Y=1207198
X3755 12270 12262 25 12296 12366 26 12380 12469 OAI221XL $T=1242000 1310770 1 0 $X=1241998 $Y=1306830
X3756 11706 12314 25 11736 11576 26 12457 12456 OAI221XL $T=1246140 1229590 1 0 $X=1246138 $Y=1225650
X3757 12270 12455 25 12172 12527 26 12538 12554 OAI221XL $T=1248440 1332910 1 0 $X=1248438 $Y=1328970
X3758 11568 12472 25 12296 12193 26 12560 12317 OAI221XL $T=1249360 1214830 0 0 $X=1249358 $Y=1214578
X3759 11706 238 25 11736 12196 26 12561 12550 OAI221XL $T=1249360 1318150 0 0 $X=1249358 $Y=1317898
X3760 12270 12459 25 11586 12196 26 12608 12616 OAI221XL $T=1251200 1325530 1 0 $X=1251198 $Y=1321590
X3761 12270 12701 25 12296 11576 26 12660 12502 OAI221XL $T=1259020 1222210 0 180 $X=1255800 $Y=1218270
X3762 12270 12634 25 11586 12641 26 12755 12853 OAI221XL $T=1258100 1318150 1 0 $X=1258098 $Y=1314210
X3763 12270 12506 25 11586 12766 26 12778 12861 OAI221XL $T=1259020 1332910 1 0 $X=1259018 $Y=1328970
X3764 12270 12821 25 12296 12914 26 12938 13068 OAI221XL $T=1266840 1288630 1 0 $X=1266838 $Y=1284690
X3765 12270 12912 25 12296 12818 26 12958 12933 OAI221XL $T=1267300 1332910 1 0 $X=1267298 $Y=1328970
X3766 11706 12856 25 11736 13033 26 13044 13067 OAI221XL $T=1271440 1244350 1 0 $X=1271438 $Y=1240410
X3767 11706 275 25 11736 12914 26 13045 13089 OAI221XL $T=1271440 1296010 1 0 $X=1271438 $Y=1292070
X3768 12270 13095 25 12296 13118 26 13128 13135 OAI221XL $T=1275580 1222210 0 0 $X=1275578 $Y=1221958
X3769 11706 12964 25 11736 13000 26 13130 13149 OAI221XL $T=1275580 1281250 0 0 $X=1275578 $Y=1280998
X3770 12270 13099 25 12296 12947 26 13132 13150 OAI221XL $T=1275580 1325530 0 0 $X=1275578 $Y=1325278
X3771 12155 13110 25 12296 13000 26 13158 13125 OAI221XL $T=1276500 1273870 1 0 $X=1276498 $Y=1269930
X3772 12270 13039 25 12296 13159 26 13172 13175 OAI221XL $T=1276960 1303390 1 0 $X=1276958 $Y=1299450
X3773 11626 282 25 11736 12947 26 13173 13187 OAI221XL $T=1276960 1325530 1 0 $X=1276958 $Y=1321590
X3774 12270 13129 25 12296 13033 26 13184 13049 OAI221XL $T=1277420 1244350 0 0 $X=1277418 $Y=1244098
X3775 12155 13097 25 12296 13079 26 13185 13115 OAI221XL $T=1277420 1259110 1 0 $X=1277418 $Y=1255170
X3776 11568 13098 25 12296 13011 26 13186 13166 OAI221XL $T=1277420 1303390 0 0 $X=1277418 $Y=1303138
X3777 11706 297 25 11736 13159 26 13234 13201 OAI221XL $T=1285240 1296010 1 180 $X=1282020 $Y=1295758
X3778 11706 13238 25 11736 13079 26 13274 13281 OAI221XL $T=1282480 1251730 0 0 $X=1282478 $Y=1251478
X3779 11706 292 25 11736 13011 26 13283 13259 OAI221XL $T=1282940 1310770 0 0 $X=1282938 $Y=1310518
X3780 12155 13258 25 12296 13228 26 13340 13004 OAI221XL $T=1285240 1266490 0 0 $X=1285238 $Y=1266238
X3781 314 12792 25 13439 312 26 13419 13299 OAI221XL $T=1293980 1185310 1 180 $X=1290760 $Y=1185058
X3782 314 13390 25 13316 312 26 13449 13375 OAI221XL $T=1296280 1273870 1 180 $X=1293060 $Y=1273618
X3783 314 12051 25 13366 312 26 13450 13365 OAI221XL $T=1296280 1310770 1 180 $X=1293060 $Y=1310518
X3784 314 12143 25 13457 312 26 13475 13645 OAI221XL $T=1293520 1222210 0 0 $X=1293518 $Y=1221958
X3785 314 13405 25 13476 312 26 13504 13564 OAI221XL $T=1294440 1244350 1 0 $X=1294438 $Y=1240410
X3786 314 12258 25 13437 312 26 13531 13555 OAI221XL $T=1295360 1347670 1 0 $X=1295358 $Y=1343730
X3787 314 12063 25 13511 312 26 13331 13469 OAI221XL $T=1298580 1185310 1 180 $X=1295360 $Y=1185058
X3788 314 12050 25 13430 312 26 13565 13253 OAI221XL $T=1302260 1281250 1 180 $X=1299040 $Y=1280998
X3789 314 12039 25 13590 312 26 13602 13652 OAI221XL $T=1299960 1229590 1 0 $X=1299958 $Y=1225650
X3790 314 13332 25 13548 312 26 13615 13627 OAI221XL $T=1299960 1251730 0 0 $X=1299958 $Y=1251478
X3791 314 12024 25 13559 312 26 13617 13647 OAI221XL $T=1299960 1332910 1 0 $X=1299958 $Y=1328970
X3792 314 12516 25 13512 312 26 13635 13614 OAI221XL $T=1300880 1200070 1 0 $X=1300878 $Y=1196130
X3793 314 12589 25 13373 312 26 13622 13692 OAI221XL $T=1302260 1185310 0 0 $X=1302258 $Y=1185058
X3794 314 12110 25 13616 312 26 13625 13612 OAI221XL $T=1305480 1318150 0 180 $X=1302260 $Y=1314210
X3795 314 12142 25 13513 312 26 13675 13673 OAI221XL $T=1303640 1214830 1 0 $X=1303638 $Y=1210890
X3796 314 12754 25 13729 312 26 13722 13672 OAI221XL $T=1315140 1200070 0 180 $X=1311920 $Y=1196130
X3797 314 13329 25 346 312 26 345 13724 OAI221XL $T=1315600 1347670 1 180 $X=1312380 $Y=1347418
X3798 8818 8931 8880 8943 25 26 8950 OA22X1 $T=1063520 1141030 1 0 $X=1063518 $Y=1137090
X3799 8954 8951 8947 8932 25 26 8930 OA22X1 $T=1066740 1177930 1 180 $X=1063980 $Y=1177678
X3800 8872 8940 8936 8946 25 26 8937 OA22X1 $T=1067200 1177930 0 180 $X=1064440 $Y=1173990
X3801 8976 9005 8980 8975 25 26 8941 OA22X1 $T=1070880 1133650 0 180 $X=1068120 $Y=1129710
X3802 8976 8936 8822 8975 25 26 9077 OA22X1 $T=1069960 1148410 1 0 $X=1069958 $Y=1144470
X3803 8947 8741 8940 8943 25 26 9120 OA22X1 $T=1069960 1148410 0 0 $X=1069958 $Y=1148158
X3804 8870 8920 8859 8931 25 26 9001 OA22X1 $T=1078240 1163170 1 180 $X=1075480 $Y=1162918
X3805 8980 9177 9243 8975 25 26 9262 OA22X1 $T=1085600 1133650 0 0 $X=1085598 $Y=1133398
X3806 8880 8741 9005 8943 25 26 9276 OA22X1 $T=1091120 1141030 0 180 $X=1088360 $Y=1137090
X3807 9531 9406 9297 9406 25 26 9218 OA22X1 $T=1097560 1207450 0 180 $X=1094800 $Y=1203510
X3808 58 9382 9686 9699 25 26 9717 OA22X1 $T=1109520 1259110 0 0 $X=1109518 $Y=1258858
X3809 38 9382 9686 9554 25 26 9745 OA22X1 $T=1109520 1281250 1 0 $X=1109518 $Y=1277310
X3810 27 9382 9686 9418 25 26 9837 OA22X1 $T=1111360 1273870 1 0 $X=1111358 $Y=1269930
X3811 63 85 9686 9782 25 26 10076 OA22X1 $T=1122860 1266490 0 0 $X=1122858 $Y=1266238
X3812 47 85 9686 10534 25 26 10535 OA22X1 $T=1149080 1266490 0 0 $X=1149078 $Y=1266238
X3813 10669 10273 85 9663 25 26 10618 OA22X1 $T=1158740 1288630 0 180 $X=1155980 $Y=1284690
X3814 10290 10791 10809 10260 25 26 10998 OA22X1 $T=1173460 1288630 0 0 $X=1173458 $Y=1288378
X3815 10888 10290 10260 10840 25 26 10974 OA22X1 $T=1182660 1281250 1 180 $X=1179900 $Y=1280998
X3816 10290 11431 11419 10260 25 26 11390 OA22X1 $T=1198760 1296010 0 180 $X=1196000 $Y=1292070
X3817 218 12005 11992 11978 25 26 11814 OA22X1 $T=1226360 1318150 1 180 $X=1223600 $Y=1317898
X3818 12039 12015 12000 11988 25 26 11842 OA22X1 $T=1226820 1236970 1 180 $X=1224060 $Y=1236718
X3819 12050 12016 12001 11989 25 26 11844 OA22X1 $T=1226820 1251730 1 180 $X=1224060 $Y=1251478
X3820 219 12016 12001 11990 25 26 11845 OA22X1 $T=1226820 1266490 0 180 $X=1224060 $Y=1262550
X3821 12051 12005 12001 11977 25 26 11813 OA22X1 $T=1226820 1288630 1 180 $X=1224060 $Y=1288378
X3822 12024 12017 12000 11991 25 26 11615 OA22X1 $T=1226820 1310770 0 180 $X=1224060 $Y=1306830
X3823 12063 12016 12001 11891 25 26 11929 OA22X1 $T=1227740 1214830 0 180 $X=1224980 $Y=1210890
X3824 12050 12015 12000 11989 25 26 11745 OA22X1 $T=1227740 1251730 0 180 $X=1224980 $Y=1247790
X3825 219 12015 12000 11990 25 26 11910 OA22X1 $T=1227740 1259110 0 180 $X=1224980 $Y=1255170
X3826 12110 12005 11992 12009 25 26 11768 OA22X1 $T=1227740 1281250 1 180 $X=1224980 $Y=1280998
X3827 12051 12017 12000 11977 25 26 11812 OA22X1 $T=1227740 1288630 0 180 $X=1224980 $Y=1284690
X3828 218 12017 12000 11978 25 26 11735 OA22X1 $T=1227740 1318150 0 180 $X=1224980 $Y=1314210
X3829 12063 12015 12000 11891 25 26 11938 OA22X1 $T=1228200 1207450 0 180 $X=1225440 $Y=1203510
X3830 12142 12016 12001 12038 25 26 11960 OA22X1 $T=1228660 1222210 0 180 $X=1225900 $Y=1218270
X3831 12110 12017 12000 12009 25 26 11746 OA22X1 $T=1230500 1273870 1 180 $X=1227740 $Y=1273618
X3832 12142 12015 12000 12038 25 26 11999 OA22X1 $T=1235100 1214830 1 180 $X=1232340 $Y=1214578
X3833 12258 12017 12000 12171 25 26 11689 OA22X1 $T=1235560 1266490 1 180 $X=1232800 $Y=1266238
X3834 12143 12015 12000 12119 25 26 11966 OA22X1 $T=1238780 1229590 1 180 $X=1236020 $Y=1229338
X3835 12258 12016 12001 12171 25 26 12115 OA22X1 $T=1238780 1273870 0 180 $X=1236020 $Y=1269930
X3836 230 12017 12000 12260 25 26 11655 OA22X1 $T=1240160 1303390 0 180 $X=1237400 $Y=1299450
X3837 228 12017 12000 12284 25 26 12271 OA22X1 $T=1241540 1318150 1 180 $X=1238780 $Y=1317898
X3838 228 12005 12117 12284 25 26 12239 OA22X1 $T=1241540 1325530 0 180 $X=1238780 $Y=1321590
X3839 230 12005 12001 12260 25 26 11972 OA22X1 $T=1245220 1303390 0 180 $X=1242460 $Y=1299450
X3840 12516 12015 12000 12323 25 26 12331 OA22X1 $T=1251200 1207450 0 180 $X=1248440 $Y=1203510
X3841 12589 12015 12000 12599 25 26 12348 OA22X1 $T=1255340 1236970 1 180 $X=1252580 $Y=1236718
X3842 252 12017 12352 12617 25 26 12538 OA22X1 $T=1255800 1332910 1 180 $X=1253040 $Y=1332658
X3843 252 12005 12117 12617 25 26 12555 OA22X1 $T=1257180 1340290 1 180 $X=1254420 $Y=1340038
X3844 12754 12016 12001 12649 25 26 12257 OA22X1 $T=1257640 1214830 0 180 $X=1254880 $Y=1210890
X3845 12754 12015 12000 12649 25 26 12560 OA22X1 $T=1260860 1207450 0 180 $X=1258100 $Y=1203510
X3846 12792 12015 12000 12726 25 26 12660 OA22X1 $T=1261320 1214830 1 180 $X=1258560 $Y=1214578
X3847 260 12017 12336 12727 25 26 12380 OA22X1 $T=1261320 1310770 0 180 $X=1258560 $Y=1306830
X3848 262 12005 12001 12728 25 26 12561 OA22X1 $T=1261320 1318150 1 180 $X=1258560 $Y=1317898
X3849 12792 12016 12001 12726 25 26 12457 OA22X1 $T=1262240 1222210 1 180 $X=1259480 $Y=1221958
X3850 260 12144 12001 12727 25 26 12718 OA22X1 $T=1262240 1303390 0 180 $X=1259480 $Y=1299450
X3851 262 12017 12336 12728 25 26 12608 OA22X1 $T=1268680 1325530 0 180 $X=1265920 $Y=1321590
X3852 285 12017 12352 13119 25 26 12778 OA22X1 $T=1279260 1332910 1 180 $X=1276500 $Y=1332658
X3853 287 12005 12117 13120 25 26 13005 OA22X1 $T=1279260 1340290 1 180 $X=1276500 $Y=1340038
X3854 296 12017 12336 13160 25 26 12755 OA22X1 $T=1280640 1318150 0 180 $X=1277880 $Y=1314210
X3855 287 12017 12352 13120 25 26 12958 OA22X1 $T=1281560 1340290 0 180 $X=1278800 $Y=1336350
X3856 299 12358 12336 13239 25 26 13186 OA22X1 $T=1284780 1303390 1 180 $X=1282020 $Y=1303138
X3857 305 12017 12336 13245 25 26 13132 OA22X1 $T=1285240 1325530 1 180 $X=1282480 $Y=1325278
X3858 305 12005 12117 13245 25 26 13173 OA22X1 $T=1286160 1325530 0 180 $X=1283400 $Y=1321590
X3859 296 12005 12117 13160 25 26 13037 OA22X1 $T=1286620 1318150 1 180 $X=1283860 $Y=1317898
X3860 13329 12144 12117 13282 25 26 13249 OA22X1 $T=1287080 1273870 0 180 $X=1284320 $Y=1269930
X3861 285 12005 12117 13119 25 26 13264 OA22X1 $T=1287080 1332910 0 180 $X=1284320 $Y=1328970
X3862 13275 301 13280 304 25 26 13331 OA22X1 $T=1284780 1192690 1 0 $X=1284778 $Y=1188750
X3863 13332 12015 12336 13292 25 26 13128 OA22X1 $T=1287540 1222210 1 180 $X=1284780 $Y=1221958
X3864 13405 12358 12336 13294 25 26 13184 OA22X1 $T=1287540 1244350 1 180 $X=1284780 $Y=1244098
X3865 313 12005 12117 13295 25 26 13130 OA22X1 $T=1287540 1281250 1 180 $X=1284780 $Y=1280998
X3866 317 12005 12117 13296 25 26 13234 OA22X1 $T=1287540 1303390 0 180 $X=1284780 $Y=1299450
X3867 13332 12144 12117 13292 25 26 13284 OA22X1 $T=1288000 1229590 1 180 $X=1285240 $Y=1229338
X3868 13390 12358 12336 13305 25 26 13185 OA22X1 $T=1288000 1259110 0 180 $X=1285240 $Y=1255170
X3869 307 12017 12336 13306 25 26 12938 OA22X1 $T=1288000 1288630 1 180 $X=1285240 $Y=1288378
X3870 307 12005 12117 13306 25 26 13045 OA22X1 $T=1288000 1296010 0 180 $X=1285240 $Y=1292070
X3871 299 12005 12117 13239 25 26 13283 OA22X1 $T=1288000 1310770 0 180 $X=1285240 $Y=1306830
X3872 13390 12144 12117 13305 25 26 13274 OA22X1 $T=1290300 1251730 0 180 $X=1287540 $Y=1247790
X3873 13405 12144 12117 13294 25 26 13044 OA22X1 $T=1290760 1244350 0 180 $X=1288000 $Y=1240410
X3874 13429 301 13458 304 25 26 13504 OA22X1 $T=1293520 1244350 0 0 $X=1293518 $Y=1244098
X3875 317 12017 12336 13296 25 26 13172 OA22X1 $T=1293520 1303390 1 0 $X=1293518 $Y=1299450
X3876 13308 301 13465 304 25 26 13419 OA22X1 $T=1296280 1192690 0 180 $X=1293520 $Y=1188750
X3877 313 12358 12336 13295 25 26 13158 OA22X1 $T=1296280 1281250 1 180 $X=1293520 $Y=1280998
X3878 13392 301 13382 304 25 26 13531 OA22X1 $T=1294440 1340290 0 0 $X=1294438 $Y=1340038
X3879 13519 301 13492 304 25 26 13450 OA22X1 $T=1297660 1318150 0 180 $X=1294900 $Y=1314210
X3880 13470 301 13491 304 25 26 13475 OA22X1 $T=1295360 1229590 1 0 $X=1295358 $Y=1225650
X3881 13329 12358 12336 13282 25 26 13340 OA22X1 $T=1295360 1266490 0 0 $X=1295358 $Y=1266238
X3882 328 301 13244 304 25 26 13449 OA22X1 $T=1298580 1281250 0 180 $X=1295820 $Y=1277310
X3883 13490 301 13510 304 25 26 13622 OA22X1 $T=1299960 1192690 1 0 $X=1299958 $Y=1188750
X3884 13568 301 13591 304 25 26 13625 OA22X1 $T=1299960 1310770 0 0 $X=1299958 $Y=1310518
X3885 13220 301 13601 304 25 26 13617 OA22X1 $T=1300420 1332910 0 0 $X=1300418 $Y=1332658
X3886 13624 301 13445 304 25 26 13565 OA22X1 $T=1303180 1288630 0 180 $X=1300420 $Y=1284690
X3887 13587 301 13600 304 25 26 13615 OA22X1 $T=1301340 1259110 1 0 $X=1301338 $Y=1255170
X3888 13649 301 13623 304 25 26 13602 OA22X1 $T=1304100 1229590 1 180 $X=1301340 $Y=1229338
X3889 13626 301 13502 304 25 26 13635 OA22X1 $T=1306860 1200070 1 0 $X=1306858 $Y=1196130
X3890 13639 301 13607 304 25 26 13722 OA22X1 $T=1310540 1200070 0 0 $X=1310538 $Y=1199818
X3891 13691 301 13663 304 25 26 13675 OA22X1 $T=1311460 1214830 0 0 $X=1311458 $Y=1214578
X3892 8835 8736 8733 25 8732 26 8679 AO22X1 $T=1044660 1177930 0 180 $X=1041900 $Y=1173990
X3893 8838 8742 8748 25 8743 26 8739 AO22X1 $T=1049260 1163170 1 180 $X=1046500 $Y=1162918
X3894 8750 8814 8734 25 8816 26 8735 AO22X1 $T=1054780 1155790 1 180 $X=1052020 $Y=1155538
X3895 9013 8749 8961 25 8952 26 8910 AO22X1 $T=1068580 1118890 0 180 $X=1065820 $Y=1114950
X3896 9013 8961 9003 25 8952 26 8970 AO22X1 $T=1071340 1118890 1 180 $X=1068580 $Y=1118638
X3897 8793 9003 9101 25 8824 26 9200 AO22X1 $T=1077320 1126270 1 0 $X=1077318 $Y=1122330
X3898 9228 8792 8935 25 9102 26 9261 AO22X1 $T=1086060 1118890 1 0 $X=1086058 $Y=1114950
X3899 9532 9542 9176 25 9573 26 9599 AO22X1 $T=1103080 1111510 0 0 $X=1103078 $Y=1111258
X3900 9532 9543 9039 25 9573 26 9564 AO22X1 $T=1103080 1118890 1 0 $X=1103078 $Y=1114950
X3901 9532 9544 9273 25 9573 26 9587 AO22X1 $T=1103080 1118890 0 0 $X=1103078 $Y=1118638
X3902 9379 9264 9555 25 8749 26 9584 AO22X1 $T=1103080 1148410 0 0 $X=1103078 $Y=1148158
X3903 9392 9625 9513 25 9363 26 9565 AO22X1 $T=1107680 1192690 0 180 $X=1104920 $Y=1188750
X3904 9532 9598 9038 25 9573 26 9696 AO22X1 $T=1105380 1104130 0 0 $X=1105378 $Y=1103878
X3905 9532 9728 9583 25 9573 26 9764 AO22X1 $T=1111820 1104130 1 0 $X=1111818 $Y=1100190
X3906 9800 9766 9756 25 9575 26 9720 AO22X1 $T=1115040 1214830 1 180 $X=1112280 $Y=1214578
X3907 9392 9774 9117 25 9363 26 9709 AO22X1 $T=1115500 1104130 1 180 $X=1112740 $Y=1103878
X3908 9532 9805 8918 25 9573 26 9838 AO22X1 $T=1115500 1096750 0 0 $X=1115498 $Y=1096498
X3909 9988 9857 9949 25 9920 26 9889 AO22X1 $T=1124700 1074610 1 180 $X=1121940 $Y=1074358
X3910 9988 9095 9968 25 9920 26 9917 AO22X1 $T=1125160 1074610 0 180 $X=1122400 $Y=1070670
X3911 9532 10024 9727 25 9573 26 10118 AO22X1 $T=1126080 1096750 0 0 $X=1126078 $Y=1096498
X3912 9988 9926 10065 25 9920 26 10079 AO22X1 $T=1127920 1059850 0 0 $X=1127918 $Y=1059598
X3913 9532 10056 9703 25 9573 26 10180 AO22X1 $T=1127920 1111510 1 0 $X=1127918 $Y=1107570
X3914 9988 9562 10105 25 9920 26 10043 AO22X1 $T=1131600 1067230 1 180 $X=1128840 $Y=1066978
X3915 9988 9900 10123 25 9920 26 10034 AO22X1 $T=1132060 1052470 1 180 $X=1129300 $Y=1052218
X3916 9988 9618 10175 25 9920 26 10150 AO22X1 $T=1134360 1052470 0 180 $X=1131600 $Y=1048530
X3917 9988 10094 10186 25 9920 26 10236 AO22X1 $T=1132520 1170550 0 0 $X=1132518 $Y=1170298
X3918 9988 9592 10210 25 9920 26 10240 AO22X1 $T=1133900 1059850 0 0 $X=1133898 $Y=1059598
X3919 9532 10267 9960 25 9573 26 10303 AO22X1 $T=1137120 1118890 1 0 $X=1137118 $Y=1114950
X3920 9392 10324 9252 25 9363 26 10283 AO22X1 $T=1141260 1170550 1 180 $X=1138500 $Y=1170298
X3921 9988 10247 10323 25 9920 26 10259 AO22X1 $T=1141720 1170550 0 180 $X=1138960 $Y=1166610
X3922 9840 9962 10471 25 10484 26 9880 AO22X1 $T=1146320 1185310 0 0 $X=1146318 $Y=1185058
X3923 9988 10433 10544 25 10484 26 10491 AO22X1 $T=1152300 1052470 1 180 $X=1149540 $Y=1052218
X3924 9988 10093 10550 25 9920 26 10527 AO22X1 $T=1152760 1059850 0 180 $X=1150000 $Y=1055910
X3925 9532 10630 9950 25 9573 26 10604 AO22X1 $T=1157820 1126270 0 180 $X=1155060 $Y=1122330
X3926 9988 10531 10636 25 10484 26 10614 AO22X1 $T=1158740 1059850 0 180 $X=1155980 $Y=1055910
X3927 9988 10762 10754 25 10484 26 10738 AO22X1 $T=1164720 1059850 0 180 $X=1161960 $Y=1055910
X3928 9988 10778 10966 25 9920 26 10802 AO22X1 $T=1175760 1052470 1 180 $X=1173000 $Y=1052218
X3929 172 11246 11217 25 166 26 165 AO22X1 $T=1188640 1332910 1 180 $X=1185880 $Y=1332658
X3930 172 11315 11325 25 166 26 178 AO22X1 $T=1190940 1332910 0 0 $X=1190938 $Y=1332658
X3931 9392 11185 11447 25 9363 26 11545 AO22X1 $T=1197840 1126270 1 0 $X=1197838 $Y=1122330
X3932 9392 11057 11452 25 9363 26 11526 AO22X1 $T=1198300 1104130 0 0 $X=1198298 $Y=1103878
X3933 9532 11144 11538 25 9363 26 11548 AO22X1 $T=1202900 1111510 0 0 $X=1202898 $Y=1111258
X3934 172 11504 11557 25 166 26 190 AO22X1 $T=1210260 1340290 1 180 $X=1207500 $Y=1340038
X3935 9392 11237 11620 25 9363 26 11726 AO22X1 $T=1207960 1111510 0 0 $X=1207958 $Y=1111258
X3936 172 11562 11619 25 166 26 198 AO22X1 $T=1208420 1340290 1 0 $X=1208418 $Y=1336350
X3937 9840 11755 11771 25 9920 26 11822 AO22X1 $T=1213940 1148410 1 0 $X=1213938 $Y=1144470
X3938 11901 11980 11561 25 11546 26 11947 AO22X1 $T=1225440 1185310 1 180 $X=1222680 $Y=1185058
X3939 9392 10923 11979 25 9363 26 12022 AO22X1 $T=1223600 1118890 1 0 $X=1223598 $Y=1114950
X3940 9392 11183 11985 25 9363 26 12065 AO22X1 $T=1224980 1104130 0 0 $X=1224978 $Y=1103878
X3941 9392 10594 12025 25 9363 26 12064 AO22X1 $T=1225440 1111510 1 0 $X=1225438 $Y=1107570
X3942 9392 10828 12026 25 9363 26 12132 AO22X1 $T=1225440 1111510 0 0 $X=1225438 $Y=1111258
X3943 9532 11058 12027 25 9363 26 12092 AO22X1 $T=1225440 1126270 1 0 $X=1225438 $Y=1122330
X3944 9532 10643 12471 25 9573 26 12517 AO22X1 $T=1247980 1096750 0 0 $X=1247978 $Y=1096498
X3945 9532 10706 12493 25 9573 26 12621 AO22X1 $T=1248440 1096750 1 0 $X=1248438 $Y=1092810
X3946 9392 10848 12513 25 9573 26 12583 AO22X1 $T=1249820 1104130 1 0 $X=1249818 $Y=1100190
X3947 9532 10742 12553 25 9573 26 12499 AO22X1 $T=1252580 1111510 0 180 $X=1249820 $Y=1107570
X3948 9532 10917 12618 25 9573 26 12648 AO22X1 $T=1253040 1118890 1 0 $X=1253038 $Y=1114950
X3949 9532 10847 12632 25 9573 26 12639 AO22X1 $T=1253960 1096750 0 0 $X=1253958 $Y=1096498
X3950 9532 10958 12633 25 9573 26 12674 AO22X1 $T=1253960 1111510 0 0 $X=1253958 $Y=1111258
X3951 298 212 295 25 290 26 13229 AO22X1 $T=1284780 1347670 1 180 $X=1282020 $Y=1347418
X3952 286 291 293 25 13256 26 13327 AO22X1 $T=1282480 1207450 1 0 $X=1282478 $Y=1203510
X3953 286 142 293 25 13257 26 13328 AO22X1 $T=1282480 1207450 0 0 $X=1282478 $Y=1207198
X3954 286 294 293 25 13273 26 13272 AO22X1 $T=1282940 1222210 1 0 $X=1282938 $Y=1218270
X3955 286 302 293 25 13314 26 13339 AO22X1 $T=1284780 1266490 1 0 $X=1284778 $Y=1262550
X3956 298 220 295 25 13315 26 13352 AO22X1 $T=1284780 1332910 0 0 $X=1284778 $Y=1332658
X3957 13247 13252 13247 25 13105 26 13326 AO22X1 $T=1288920 1170550 0 0 $X=1288918 $Y=1170298
X3958 286 153 293 25 13379 26 13348 AO22X1 $T=1291680 1222210 0 180 $X=1288920 $Y=1218270
X3959 286 151 293 25 13093 26 13503 AO22X1 $T=1291220 1200070 0 0 $X=1291218 $Y=1199818
X3960 286 311 293 25 13505 26 13364 AO22X1 $T=1294900 1259110 0 0 $X=1294898 $Y=1258858
X3961 298 326 295 25 13260 26 13514 AO22X1 $T=1294900 1325530 1 0 $X=1294898 $Y=1321590
X3962 286 187 293 25 13380 26 13313 AO22X1 $T=1298580 1236970 1 180 $X=1295820 $Y=1236718
X3963 286 161 293 25 13608 26 13644 AO22X1 $T=1299960 1207450 1 0 $X=1299958 $Y=1203510
X3964 298 211 295 25 13603 26 13653 AO22X1 $T=1301340 1325530 1 0 $X=1301338 $Y=1321590
X3965 286 333 295 25 13351 26 13585 AO22X1 $T=1304100 1303390 0 180 $X=1301340 $Y=1299450
X3966 286 182 293 25 13338 26 13530 AO22X1 $T=1302260 1244350 0 0 $X=1302258 $Y=1244098
X3967 8836 26 8679 8739 8735 25 8825 NOR4X1 $T=1045580 1170550 0 180 $X=1043280 $Y=1166610
X3968 8869 26 8879 8905 8910 25 8966 NOR4X1 $T=1060300 1118890 0 0 $X=1060298 $Y=1118638
X3969 9066 26 8971 9004 8970 25 9086 NOR4X1 $T=1071340 1126270 1 180 $X=1069040 $Y=1126018
X3970 9533 26 9539 9229 9564 25 9679 NOR4X1 $T=1103080 1155790 0 0 $X=1103078 $Y=1155538
X3971 9364 26 9545 9556 9565 25 9697 NOR4X1 $T=1103080 1185310 1 0 $X=1103078 $Y=1181370
X3972 9769 26 9492 9145 9696 25 9799 NOR4X1 $T=1112740 1155790 1 180 $X=1110440 $Y=1155538
X3973 10199 26 105 106 10302 25 10363 NOR4X1 $T=1138040 1347670 0 0 $X=1138038 $Y=1347418
X3974 9559 26 25 9375 9350 9394 NAND3BX1 $T=1097560 1244350 0 180 $X=1095260 $Y=1240410
X3975 9668 26 25 9687 9700 9375 NAND3BX1 $T=1109520 1303390 1 0 $X=1109518 $Y=1299450
X3976 44 26 25 9375 9438 9667 NAND3BX1 $T=1111820 1229590 1 180 $X=1109520 $Y=1229338
X3977 9720 26 25 9698 9546 9660 NAND3BX1 $T=1112280 1222210 1 180 $X=1109980 $Y=1221958
X3978 8868 8904 8918 25 26 XOR2X1 $T=1060300 1096750 1 0 $X=1060298 $Y=1092810
X3979 8979 9084 9117 25 26 XOR2X1 $T=1075940 1089370 0 0 $X=1075938 $Y=1089118
X3980 9140 9115 9095 25 26 XOR2X1 $T=1079160 1067230 0 180 $X=1075940 $Y=1063290
X3981 9255 9246 9291 25 26 XOR2X1 $T=1087440 1111510 1 0 $X=1087438 $Y=1107570
X3982 9342 9469 9513 25 26 XOR2X1 $T=1099860 1192690 1 0 $X=1099858 $Y=1188750
X3983 9474 9581 9618 25 26 XOR2X1 $T=1104460 1052470 0 0 $X=1104458 $Y=1052218
X3984 9586 9657 9727 25 26 XOR2X1 $T=1110440 1096750 1 0 $X=1110438 $Y=1092810
X3985 9547 9723 9691 25 26 XOR2X1 $T=1113660 1296010 1 180 $X=1110440 $Y=1295758
X3986 9850 9826 9766 25 26 XOR2X1 $T=1118720 1222210 0 180 $X=1115500 $Y=1218270
X3987 9905 9894 9950 25 26 XOR2X1 $T=1121480 1096750 1 0 $X=1121478 $Y=1092810
X3988 10856 10798 10778 25 26 XOR2X1 $T=1166560 1037710 0 180 $X=1163340 $Y=1033770
X3989 11432 11595 11619 25 26 XOR2X1 $T=1206120 1332910 0 0 $X=1206118 $Y=1332658
X3990 11687 11614 11447 25 26 XOR2X1 $T=1209340 1126270 0 180 $X=1206120 $Y=1122330
X3991 12181 12166 12027 25 26 XOR2X1 $T=1234640 1126270 0 180 $X=1231420 $Y=1122330
X3992 12241 12180 12025 25 26 XOR2X1 $T=1235560 1052470 1 180 $X=1232340 $Y=1052218
X3993 12616 12550 12530 25 26 XOR2X1 $T=1252580 1318150 0 180 $X=1249360 $Y=1314210
X3994 12684 12715 12618 25 26 XOR2X1 $T=1258100 1074610 0 0 $X=1258098 $Y=1074358
X3995 12708 12743 12553 25 26 XOR2X1 $T=1259020 1104130 0 0 $X=1259018 $Y=1103878
X3996 12932 12853 12871 25 26 XOR2X1 $T=1269140 1318150 0 180 $X=1265920 $Y=1314210
X3997 13089 13068 13126 25 26 XOR2X1 $T=1275580 1288630 1 0 $X=1275578 $Y=1284690
X3998 13517 13489 12563 25 26 XOR2X1 $T=1297660 1133650 0 180 $X=1294440 $Y=1129710
X3999 13681 13709 12919 25 26 XOR2X1 $T=1310080 1111510 1 0 $X=1310078 $Y=1107570
X4000 8837 8745 25 8862 26 8878 OAI21XL $T=1058920 1104130 1 0 $X=1058918 $Y=1100190
X4001 9008 8903 25 8939 26 8977 OAI21XL $T=1070880 1081990 0 180 $X=1069040 $Y=1078050
X4002 8945 9042 25 8837 26 8972 OAI21XL $T=1072260 1104130 0 180 $X=1070420 $Y=1100190
X4003 8969 9010 25 9123 26 9239 OAI21XL $T=1077320 1214830 1 0 $X=1077318 $Y=1210890
X4004 9210 9085 25 9106 26 9092 OAI21XL $T=1079620 1104130 1 180 $X=1077780 $Y=1103878
X4005 9219 9220 25 9088 26 9100 OAI21XL $T=1085140 1089370 1 180 $X=1083300 $Y=1089118
X4006 9357 9249 25 9241 26 9139 OAI21XL $T=1087900 1067230 1 180 $X=1086060 $Y=1066978
X4007 9231 9250 25 9236 26 9260 OAI21XL $T=1086520 1081990 1 0 $X=1086518 $Y=1078050
X4008 9153 9255 25 9210 26 9216 OAI21XL $T=1088360 1104130 1 180 $X=1086520 $Y=1103878
X4009 9300 9342 25 9332 26 9237 OAI21XL $T=1094340 1192690 0 180 $X=1092500 $Y=1188750
X4010 9440 9362 25 9339 26 9118 OAI21XL $T=1095260 1104130 0 180 $X=1093420 $Y=1100190
X4011 9352 9471 25 9357 26 9485 OAI21XL $T=1098940 1067230 1 0 $X=1098938 $Y=1063290
X4012 9359 9335 25 9394 26 9540 OAI21XL $T=1098940 1214830 0 0 $X=1098938 $Y=1214578
X4013 9355 9299 25 9440 26 9486 OAI21XL $T=1099400 1096750 0 0 $X=1099398 $Y=1096498
X4014 9326 9480 25 9333 26 9503 OAI21XL $T=1099400 1214830 1 0 $X=1099398 $Y=1210890
X4015 9516 9475 25 9476 26 9347 OAI21XL $T=1101240 1081990 0 180 $X=1099400 $Y=1078050
X4016 9401 9105 25 9501 26 9530 OAI21XL $T=1100320 1052470 0 0 $X=1100318 $Y=1052218
X4017 9505 9586 25 9516 26 9615 OAI21XL $T=1104920 1089370 1 0 $X=1104918 $Y=1085430
X4018 9621 9596 25 9582 26 9577 OAI21XL $T=1106760 1067230 0 180 $X=1104920 $Y=1063290
X4019 9715 9714 25 9677 26 9568 OAI21XL $T=1112740 1045090 0 180 $X=1110900 $Y=1041150
X4020 9668 9821 25 9687 26 9739 OAI21XL $T=1117800 1303390 0 180 $X=1115960 $Y=1299450
X4021 9835 9784 25 9818 26 9707 OAI21XL $T=1118260 1059850 1 180 $X=1116420 $Y=1059598
X4022 9752 9849 25 9835 26 9865 OAI21XL $T=1117800 1052470 1 0 $X=1117798 $Y=1048530
X4023 9688 9819 25 9621 26 9898 OAI21XL $T=1121020 1067230 0 0 $X=1121018 $Y=1066978
X4024 9978 9785 25 9820 26 9373 OAI21XL $T=1122860 1081990 1 180 $X=1121020 $Y=1081738
X4025 10073 10140 25 10109 26 9899 OAI21XL $T=1132060 1200070 1 180 $X=1130220 $Y=1199818
X4026 102 10103 25 110 26 10293 OAI21XL $T=1136660 1340290 1 0 $X=1136658 $Y=1336350
X4027 103 9595 25 110 26 10320 OAI21XL $T=1138040 1310770 0 0 $X=1138038 $Y=1310518
X4028 10392 10294 25 10276 26 10179 OAI21XL $T=1139880 1045090 1 180 $X=1138040 $Y=1044838
X4029 103 10054 25 110 26 10256 OAI21XL $T=1142180 1332910 0 180 $X=1140340 $Y=1328970
X4030 103 10041 25 110 26 10249 OAI21XL $T=1140800 1332910 0 0 $X=1140798 $Y=1332658
X4031 103 10422 25 110 26 10440 OAI21XL $T=1144480 1303390 0 0 $X=1144478 $Y=1303138
X4032 103 10424 25 110 26 10437 OAI21XL $T=1144480 1318150 0 0 $X=1144478 $Y=1317898
X4033 10336 10429 25 10392 26 10405 OAI21XL $T=1146320 1045090 1 180 $X=1144480 $Y=1044838
X4034 103 10157 25 110 26 10335 OAI21XL $T=1145400 1325530 1 0 $X=1145398 $Y=1321590
X4035 103 10271 25 110 26 10488 OAI21XL $T=1146780 1340290 1 0 $X=1146778 $Y=1336350
X4036 103 10515 25 110 26 10589 OAI21XL $T=1148620 1303390 0 0 $X=1148618 $Y=1303138
X4037 103 10301 25 110 26 10149 OAI21XL $T=1151380 1325530 1 0 $X=1151378 $Y=1321590
X4038 10583 10573 25 10564 26 10200 OAI21XL $T=1153680 1037710 1 180 $X=1151840 $Y=1037458
X4039 103 10446 25 110 26 120 OAI21XL $T=1155520 1340290 1 0 $X=1155518 $Y=1336350
X4040 103 10655 25 110 26 10522 OAI21XL $T=1159200 1325530 0 180 $X=1157360 $Y=1321590
X4041 103 10581 25 110 26 10736 OAI21XL $T=1161040 1318150 1 0 $X=1161038 $Y=1314210
X4042 103 10582 25 110 26 10737 OAI21XL $T=1164720 1332910 1 180 $X=1162880 $Y=1332658
X4043 103 10722 25 110 26 10801 OAI21XL $T=1163800 1318150 1 0 $X=1163798 $Y=1314210
X4044 103 10795 25 110 26 10842 OAI21XL $T=1164260 1310770 1 0 $X=1164258 $Y=1306830
X4045 146 10983 25 11053 26 11011 OAI21XL $T=1174840 1340290 0 0 $X=1174838 $Y=1340038
X4046 11385 11422 25 11433 26 11397 OAI21XL $T=1196920 1325530 1 0 $X=1196918 $Y=1321590
X4047 11456 11150 25 11580 26 11606 OAI21XL $T=1207040 1347670 1 0 $X=1207038 $Y=1343730
X4048 11732 11616 25 11601 26 11567 OAI21XL $T=1208880 1104130 1 180 $X=1207040 $Y=1103878
X4049 11601 11749 25 11765 26 11776 OAI21XL $T=1213940 1104130 0 0 $X=1213938 $Y=1103878
X4050 202 11786 25 11770 26 11754 OAI21XL $T=1216240 1347670 1 180 $X=1214400 $Y=1347418
X4051 11614 11798 25 11839 26 11764 OAI21XL $T=1215320 1118890 1 0 $X=1215318 $Y=1114950
X4052 11862 11984 25 11799 26 12008 OAI21XL $T=1224520 1177930 0 0 $X=1224518 $Y=1177678
X4053 12223 12035 25 12141 26 12122 OAI21XL $T=1233720 1104130 1 180 $X=1231880 $Y=1103878
X4054 11828 11437 25 12134 26 12183 OAI21XL $T=1232800 1177930 0 0 $X=1232798 $Y=1177678
X4055 12219 12077 25 12182 26 12312 OAI21XL $T=1239240 1163170 0 0 $X=1239238 $Y=1162918
X4056 12236 12266 25 12307 26 12209 OAI21XL $T=1242920 1111510 1 180 $X=1241080 $Y=1111258
X4057 12302 11809 25 12377 26 12381 OAI21XL $T=1243380 1089370 0 0 $X=1243378 $Y=1089118
X4058 12141 12333 25 12363 26 12342 OAI21XL $T=1245220 1104130 0 180 $X=1243380 $Y=1100190
X4059 12460 12466 25 12600 26 12350 OAI21XL $T=1248900 1067230 1 0 $X=1248898 $Y=1063290
X4060 12182 12249 25 12391 26 12547 OAI21XL $T=1249820 1163170 0 0 $X=1249818 $Y=1162918
X4061 12551 12552 25 12535 26 12355 OAI21XL $T=1252120 1081990 0 180 $X=1250280 $Y=1078050
X4062 12545 12704 25 12714 26 12671 OAI21XL $T=1260400 1052470 1 180 $X=1258560 $Y=1052218
X4063 12763 12546 25 12716 26 12707 OAI21XL $T=1260400 1081990 1 180 $X=1258560 $Y=1081738
X4064 12539 12546 25 12552 26 12454 OAI21XL $T=1260860 1081990 0 180 $X=1259020 $Y=1078050
X4065 12604 12762 25 12750 26 12650 OAI21XL $T=1261780 1067230 0 180 $X=1259940 $Y=1063290
X4066 12691 12546 25 12673 26 12742 OAI21XL $T=1262240 1089370 1 180 $X=1260400 $Y=1089118
X4067 12673 12880 25 12982 26 13003 OAI21XL $T=1271440 1089370 1 0 $X=1271438 $Y=1085430
X4068 12881 13058 25 13100 26 13013 OAI21XL $T=1277880 1096750 1 180 $X=1276040 $Y=1096498
X4069 13104 13054 25 12868 26 13216 OAI21XL $T=1277420 1059850 0 0 $X=1277418 $Y=1059598
X4070 13261 13251 25 13232 26 13236 OAI21XL $T=1284780 1067230 1 180 $X=1282940 $Y=1066978
X4071 12815 11295 25 13304 26 13252 OAI21XL $T=1283860 1163170 1 0 $X=1283858 $Y=1159230
X4072 13372 13431 25 13361 26 13309 OAI21XL $T=1292600 1089370 0 180 $X=1290760 $Y=1085430
X4073 13440 13477 25 13486 26 13553 OAI21XL $T=1295360 1067230 1 0 $X=1295358 $Y=1063290
X4074 13474 13448 25 13488 26 13597 OAI21XL $T=1299500 1118890 1 0 $X=1299498 $Y=1114950
X4075 13619 12700 25 13596 26 13532 OAI21XL $T=1302720 1111510 1 180 $X=1300880 $Y=1111258
X4076 13562 13501 25 13427 26 13621 OAI21XL $T=1301340 1133650 0 0 $X=1301338 $Y=1133398
X4077 13446 13431 25 13477 26 13595 OAI21XL $T=1305020 1081990 1 180 $X=1303180 $Y=1081738
X4078 13418 13506 25 13459 26 13620 OAI21XL $T=1305020 1104130 0 180 $X=1303180 $Y=1100190
X4079 13582 13681 25 13474 26 13581 OAI21XL $T=1307320 1111510 1 180 $X=1305480 $Y=1111258
X4080 13711 13431 25 13714 26 13737 OAI21XL $T=1311000 1089370 1 0 $X=1310998 $Y=1085430
X4081 11389 11739 11627 25 26 11795 MX2X1 $T=1213480 1081990 0 0 $X=1213478 $Y=1081738
X4082 11389 11940 11738 25 26 11892 MX2X1 $T=1223140 1059850 0 180 $X=1219460 $Y=1055910
X4083 11389 12151 11958 25 26 12040 MX2X1 $T=1233720 1037710 0 180 $X=1230040 $Y=1033770
X4084 16519 607 16530 25 26 13971 MX2X1 $T=1582400 1288630 0 180 $X=1578720 $Y=1284690
X4085 16519 16544 16551 25 26 13919 MX2X1 $T=1582860 1288630 1 180 $X=1579180 $Y=1288378
X4086 603 613 16586 25 26 355 MX2X1 $T=1590680 1340290 0 180 $X=1587000 $Y=1336350
X4087 16519 16724 16710 25 26 13739 MX2X1 $T=1604940 1236970 1 180 $X=1601260 $Y=1236718
X4088 52 9419 9566 25 26 XOR2XL $T=1102620 1332910 1 0 $X=1102618 $Y=1328970
X4089 59 31 9536 25 26 XOR2XL $T=1105840 1332910 1 180 $X=1102620 $Y=1332658
X4090 60 31 9724 25 26 XOR2XL $T=1109980 1347670 1 0 $X=1109978 $Y=1343730
X4091 9819 9810 9857 25 26 XOR2XL $T=1116880 1074610 1 0 $X=1116878 $Y=1070670
X4092 78 9419 9860 25 26 XOR2XL $T=1116880 1332910 0 0 $X=1116878 $Y=1332658
X4093 69 53 10199 25 26 XOR2XL $T=1132520 1347670 1 0 $X=1132518 $Y=1343730
X4094 10140 10218 10247 25 26 XOR2XL $T=1134820 1192690 0 0 $X=1134818 $Y=1192438
X4095 71 59 10302 25 26 XOR2XL $T=1141720 1347670 0 180 $X=1138500 $Y=1343730
X4096 68 52 10455 25 26 XOR2XL $T=1144480 1340290 0 0 $X=1144478 $Y=1340038
X4097 10429 10483 10531 25 26 XOR2XL $T=1148620 1045090 1 0 $X=1148618 $Y=1041150
X4098 11616 11630 11452 25 26 XOR2XL $T=1209800 1104130 0 180 $X=1206580 $Y=1100190
X4099 11869 11862 11755 25 26 XOR2XL $T=1218540 1177930 1 180 $X=1215320 $Y=1177678
X4100 12035 12006 11985 25 26 XOR2XL $T=1226820 1096750 1 180 $X=1223600 $Y=1096498
X4101 12077 12049 11849 25 26 XOR2XL $T=1228200 1170550 0 180 $X=1224980 $Y=1166610
X4102 12546 12536 12513 25 26 XOR2XL $T=1251660 1089370 1 180 $X=1248440 $Y=1089118
X4103 12466 12511 12471 25 26 XOR2XL $T=1249360 1074610 0 0 $X=1249358 $Y=1074358
X4104 13718 13468 13163 25 26 XOR2XL $T=1296280 1081990 0 180 $X=1293060 $Y=1078050
X4105 13431 13464 13121 25 26 XOR2XL $T=1294440 1081990 0 0 $X=1294438 $Y=1081738
X4106 8734 8742 26 8732 8750 8737 8748 8747 25 AOI222XL $T=1046960 1133650 1 0 $X=1046958 $Y=1129710
X4107 8824 8816 26 8814 8793 8792 8749 8746 25 AOI222XL $T=1052020 1118890 1 180 $X=1048340 $Y=1118638
X4108 8838 8871 26 8883 8911 8743 8736 8744 25 AOI222XL $T=1059840 1163170 1 0 $X=1059838 $Y=1159230
X4109 8748 8750 26 8743 8742 8814 8734 8933 25 AOI222XL $T=1063980 1155790 1 0 $X=1063978 $Y=1151850
X4110 9003 9013 26 8961 8935 8952 9101 8857 25 AOI222XL $T=1074560 1118890 0 0 $X=1074558 $Y=1118638
X4111 8814 9013 26 8748 8935 8952 8816 9089 25 AOI222XL $T=1076400 1118890 1 0 $X=1076398 $Y=1114950
X4112 9228 9013 26 9101 8935 8952 9102 8938 25 AOI222XL $T=1080540 1126270 1 180 $X=1076860 $Y=1126018
X4113 9102 9013 26 9228 8935 8952 9270 9256 25 AOI222XL $T=1085600 1126270 0 0 $X=1085598 $Y=1126018
X4114 8871 8824 26 9257 8883 8736 8792 9468 25 AOI222XL $T=1094340 1141030 1 0 $X=1094338 $Y=1137090
X4115 9194 9237 9137 25 26 9147 AO21X1 $T=1081460 1192690 1 180 $X=1079160 $Y=1192438
X4116 9344 9074 9360 25 26 9435 AO21X1 $T=1093420 1222210 1 0 $X=1093418 $Y=1218270
X4117 9487 9429 8980 25 26 9387 AO21X1 $T=1098480 1126270 1 180 $X=1096180 $Y=1126018
X4118 9487 9685 9005 25 26 9478 AO21X1 $T=1106760 1133650 0 180 $X=1104460 $Y=1129710
X4119 11245 168 11334 25 26 11293 AO21X1 $T=1191400 1325530 0 0 $X=1191398 $Y=1325278
X4120 11564 168 11606 25 26 193 AO21X1 $T=1206580 1347670 0 0 $X=1206578 $Y=1347418
X4121 13047 13108 13107 25 26 13012 AO21X1 $T=1278340 1052470 1 180 $X=1276040 $Y=1052218
X4122 13708 13737 13715 25 26 13520 AO21X1 $T=1313760 1096750 1 180 $X=1311460 $Y=1096498
X4123 9352 9357 25 26 9391 NAND2BXL $T=1094800 1067230 0 0 $X=1094798 $Y=1066978
X4124 9270 9806 25 26 9886 NAND2BXL $T=1115500 1200070 1 0 $X=1115498 $Y=1196130
X4125 10336 10392 25 26 10483 NAND2BXL $T=1144480 1045090 1 0 $X=1144478 $Y=1041150
X4126 11147 11926 25 26 12134 NAND2BXL $T=1232800 1185310 1 0 $X=1232798 $Y=1181370
X4127 11243 12943 25 26 13174 NAND2BXL $T=1284320 1177930 0 180 $X=1282480 $Y=1173990
X4128 11087 12857 25 26 13325 NAND2BXL $T=1283400 1155790 1 0 $X=1283398 $Y=1151850
X4129 11244 12929 25 26 13304 NAND2BXL $T=1295360 1163170 1 0 $X=1295358 $Y=1159230
X4130 9087 9069 9104 30 32 9202 34 26 25 SDFFRX2 $T=1074560 1325530 0 0 $X=1074558 $Y=1325278
X4131 9298 9069 9274 30 32 9104 31 26 25 SDFFRX2 $T=1091580 1332910 0 180 $X=1079160 $Y=1328970
X4132 9170 8732 25 9122 26 9108 9010 OAI211X1 $T=1079620 1214830 1 180 $X=1077320 $Y=1214578
X4133 11980 11901 25 11995 26 11947 12184 OAI211X1 $T=1235560 1185310 1 180 $X=1233260 $Y=1185058
X4134 13065 11344 25 13165 26 13174 12753 OAI211X1 $T=1277420 1177930 1 0 $X=1277418 $Y=1173990
X4135 12941 11225 25 13353 26 13325 13248 OAI211X1 $T=1289840 1148410 0 180 $X=1287540 $Y=1144470
X4136 10122 9802 10067 26 10044 10040 25 AOI2BB2X1 $T=1129760 1244350 1 180 $X=1127000 $Y=1244098
X4137 10147 9782 10067 26 10033 10077 25 AOI2BB2X1 $T=1131600 1273870 1 180 $X=1128840 $Y=1273618
X4138 9953 9915 10141 26 10081 9914 25 AOI2BB2X1 $T=1132060 1310770 1 180 $X=1129300 $Y=1310518
X4139 10147 9553 10067 26 10035 10239 25 AOI2BB2X1 $T=1132980 1266490 1 0 $X=1132978 $Y=1262550
X4140 10147 9418 10067 26 10126 10280 25 AOI2BB2X1 $T=1136660 1273870 0 0 $X=1136658 $Y=1273618
X4141 10147 9554 10067 26 10082 10396 25 AOI2BB2X1 $T=1137120 1281250 0 0 $X=1137118 $Y=1280998
X4142 10122 10003 10067 26 10311 10326 25 AOI2BB2X1 $T=1138040 1236970 0 0 $X=1138038 $Y=1236718
X4143 10147 9699 10067 26 10354 10541 25 AOI2BB2X1 $T=1144940 1266490 1 0 $X=1144938 $Y=1262550
X4144 10122 10408 10067 26 10415 10419 25 AOI2BB2X1 $T=1150460 1214830 0 180 $X=1147700 $Y=1210890
X4145 10122 10300 10067 26 10487 10570 25 AOI2BB2X1 $T=1151380 1214830 0 0 $X=1151378 $Y=1214578
X4146 10122 10539 10067 26 10596 10639 25 AOI2BB2X1 $T=1153220 1229590 1 0 $X=1153218 $Y=1225650
X4147 10147 10534 10067 26 10430 10621 25 AOI2BB2X1 $T=1154600 1281250 0 0 $X=1154598 $Y=1280998
X4148 10122 9974 10067 26 10568 10749 25 AOI2BB2X1 $T=1155060 1244350 1 0 $X=1155058 $Y=1240410
X4149 10122 10420 10067 26 10567 10721 25 AOI2BB2X1 $T=1157820 1251730 1 0 $X=1157818 $Y=1247790
X4150 10122 10703 10067 26 10705 10654 25 AOI2BB2X1 $T=1164260 1214830 0 180 $X=1161500 $Y=1210890
X4151 10122 10704 10067 26 10985 10964 25 AOI2BB2X1 $T=1173460 1207450 0 0 $X=1173458 $Y=1207198
X4152 10122 11091 10067 26 10824 11069 25 AOI2BB2X1 $T=1181280 1207450 1 180 $X=1178520 $Y=1207198
X4153 8913 8974 9038 26 25 XNOR2X1 $T=1069500 1104130 0 0 $X=1069498 $Y=1103878
X4154 8972 8962 9039 26 25 XNOR2X1 $T=1069500 1111510 0 0 $X=1069498 $Y=1111258
X4155 9147 9082 9074 26 25 XNOR2X1 $T=1077780 1222210 1 180 $X=1074560 $Y=1221958
X4156 9216 9154 9176 26 25 XNOR2X1 $T=1083300 1111510 0 180 $X=1080080 $Y=1107570
X4157 9237 9224 9273 26 25 XNOR2X1 $T=1086520 1192690 1 0 $X=1086518 $Y=1188750
X4158 9260 9266 9252 26 25 XNOR2X1 $T=1089740 1177930 1 180 $X=1086520 $Y=1177678
X4159 9486 9397 9374 26 25 XNOR2X1 $T=1097560 1111510 1 180 $X=1094340 $Y=1111258
X4160 9485 9414 9562 26 25 XNOR2X1 $T=1102620 1067230 0 0 $X=1102618 $Y=1066978
X4161 9281 9517 9583 26 25 XNOR2X1 $T=1103540 1104130 1 0 $X=1103538 $Y=1100190
X4162 9615 9661 9703 26 25 XNOR2X1 $T=1109520 1089370 0 0 $X=1109518 $Y=1089118
X4163 9865 9887 9900 26 25 XNOR2X1 $T=1119640 1052470 0 0 $X=1119638 $Y=1052218
X4164 9898 9883 9926 26 25 XNOR2X1 $T=1121020 1067230 1 0 $X=1121018 $Y=1063290
X4165 9199 9933 9960 26 25 XNOR2X1 $T=1121940 1089370 0 0 $X=1121938 $Y=1089118
X4166 10405 10277 10433 26 25 XNOR2X1 $T=1144020 1052470 0 0 $X=1144018 $Y=1052218
X4167 11293 11131 11217 26 25 XNOR2X1 $T=1188640 1332910 0 180 $X=1185420 $Y=1328970
X4168 11343 11523 11557 26 25 XNOR2X1 $T=1202900 1340290 1 0 $X=1202898 $Y=1336350
X4169 11567 11609 11620 26 25 XNOR2X1 $T=1206580 1111510 1 0 $X=1206578 $Y=1107570
X4170 11767 11623 11602 26 25 XNOR2X1 $T=1209800 1273870 0 180 $X=1206580 $Y=1269930
X4171 11647 11624 11603 26 25 XNOR2X1 $T=1209800 1303390 1 180 $X=1206580 $Y=1303138
X4172 11787 11758 11723 26 25 XNOR2X1 $T=1215780 1288630 1 180 $X=1212560 $Y=1288378
X4173 11830 11793 11730 26 25 XNOR2X1 $T=1217160 1318150 0 180 $X=1213940 $Y=1314210
X4174 11864 11769 11748 26 25 XNOR2X1 $T=1218080 1303390 0 180 $X=1214860 $Y=1299450
X4175 11784 11757 11801 26 25 XNOR2X1 $T=1215320 1273870 1 0 $X=1215318 $Y=1269930
X4176 11872 11843 11897 26 25 XNOR2X1 $T=1218540 1251730 1 0 $X=1218538 $Y=1247790
X4177 11893 11904 11920 26 25 XNOR2X1 $T=1219460 1244350 1 0 $X=1219458 $Y=1240410
X4178 11873 11906 11829 26 25 XNOR2X1 $T=1219460 1259110 0 0 $X=1219458 $Y=1258858
X4179 11802 11971 11986 26 25 XNOR2X1 $T=1223140 1207450 0 0 $X=1223138 $Y=1207198
X4180 11803 11959 11987 26 25 XNOR2X1 $T=1223140 1229590 0 0 $X=1223138 $Y=1229338
X4181 11919 11981 11982 26 25 XNOR2X1 $T=1223600 1222210 0 0 $X=1223598 $Y=1221958
X4182 12122 12145 12026 26 25 XNOR2X1 $T=1231420 1111510 1 0 $X=1231418 $Y=1107570
X4183 12312 12298 12268 26 25 XNOR2X1 $T=1241540 1163170 0 180 $X=1238320 $Y=1159230
X4184 12294 12317 12332 26 25 XNOR2X1 $T=1240160 1222210 1 0 $X=1240158 $Y=1218270
X4185 12305 12324 12343 26 25 XNOR2X1 $T=1240620 1214830 0 0 $X=1240618 $Y=1214578
X4186 12245 12346 12356 26 25 XNOR2X1 $T=1241540 1244350 1 0 $X=1241538 $Y=1240410
X4187 12456 12502 12351 26 25 XNOR2X1 $T=1248440 1222210 0 0 $X=1248438 $Y=1221958
X4188 12246 12470 12526 26 25 XNOR2X1 $T=1248440 1310770 0 0 $X=1248438 $Y=1310518
X4189 12350 12528 12493 26 25 XNOR2X1 $T=1251660 1059850 1 180 $X=1248440 $Y=1059598
X4190 12504 12469 12549 26 25 XNOR2X1 $T=1249360 1310770 1 0 $X=1249358 $Y=1306830
X4191 12519 12554 12662 26 25 XNOR2X1 $T=1254420 1325530 0 0 $X=1254418 $Y=1325278
X4192 12742 12663 12633 26 25 XNOR2X1 $T=1257640 1096750 0 180 $X=1254420 $Y=1092810
X4193 12707 12756 12632 26 25 XNOR2X1 $T=1259480 1096750 0 0 $X=1259478 $Y=1096498
X4194 12883 12861 12848 26 25 XNOR2X1 $T=1267300 1332910 1 180 $X=1264080 $Y=1332658
X4195 13012 12910 12873 26 25 XNOR2X1 $T=1269140 1052470 0 180 $X=1265920 $Y=1048530
X4196 12995 12933 12879 26 25 XNOR2X1 $T=1270060 1325530 1 180 $X=1266840 $Y=1325278
X4197 13016 13004 12984 26 25 XNOR2X1 $T=1272820 1266490 1 180 $X=1269600 $Y=1266238
X4198 13108 13035 12940 26 25 XNOR2X1 $T=1274660 1059850 0 180 $X=1271440 $Y=1055910
X4199 13067 13049 13021 26 25 XNOR2X1 $T=1275120 1244350 1 180 $X=1271900 $Y=1244098
X4200 13281 13115 13096 26 25 XNOR2X1 $T=1278340 1251730 0 180 $X=1275120 $Y=1247790
X4201 13149 13125 13103 26 25 XNOR2X1 $T=1278800 1281250 0 180 $X=1275580 $Y=1277310
X4202 13243 13146 13036 26 25 XNOR2X1 $T=1279720 1074610 0 180 $X=1276500 $Y=1070670
X4203 13187 13150 13001 26 25 XNOR2X1 $T=1279720 1318150 1 180 $X=1276500 $Y=1317898
X4204 13038 13135 13124 26 25 XNOR2X1 $T=1276960 1229590 1 0 $X=1276958 $Y=1225650
X4205 13259 13166 13131 26 25 XNOR2X1 $T=1280180 1310770 0 180 $X=1276960 $Y=1306830
X4206 13201 13175 13136 26 25 XNOR2X1 $T=1280640 1296010 1 180 $X=1277420 $Y=1295758
X4207 13309 13279 13164 26 25 XNOR2X1 $T=1286620 1089370 0 180 $X=1283400 $Y=1085430
X4208 13520 13487 13122 26 25 XNOR2X1 $T=1297660 1096750 1 180 $X=1294440 $Y=1096498
X4209 13581 13493 12794 26 25 XNOR2X1 $T=1297660 1111510 1 180 $X=1294440 $Y=1111258
X4210 13737 13730 13022 26 25 XNOR2X1 $T=1314680 1096750 0 180 $X=1311460 $Y=1092810
X4211 9536 26 9558 25 9566 9585 NOR3X1 $T=1103080 1340290 0 0 $X=1103078 $Y=1340038
X4212 9724 26 9558 25 9860 84 NOR3X1 $T=1116420 1347670 1 0 $X=1116418 $Y=1343730
X4213 9196 26 10469 25 10470 9334 NOR3X1 $T=1146780 1170550 1 0 $X=1146778 $Y=1166610
X4214 10486 26 10469 25 9196 9169 NOR3X1 $T=1148620 1170550 1 180 $X=1146780 $Y=1170298
X4215 10530 26 10470 25 9196 9043 NOR3X1 $T=1148620 1177930 0 180 $X=1146780 $Y=1173990
X4216 10486 26 9196 25 10530 9132 NOR3X1 $T=1148620 1177930 0 0 $X=1148618 $Y=1177678
X4217 9138 9005 8982 25 26 9081 AO21XL $T=1078240 1200070 1 180 $X=1075940 $Y=1199818
X4218 44 31 42 25 26 9298 AO21XL $T=1096640 1332910 1 180 $X=1094340 $Y=1332658
X4219 74 112 10166 25 26 10141 AO21XL $T=1139880 1318150 0 180 $X=1137580 $Y=1314210
X4220 13463 13595 13473 25 26 13243 AO21XL $T=1297200 1074610 0 180 $X=1294900 $Y=1070670
X4221 8863 8878 26 8877 25 8903 AOI21X1 $T=1062600 1081990 0 180 $X=1060300 $Y=1078050
X4222 8923 8913 26 8878 25 8868 AOI21X1 $T=1062600 1096750 1 180 $X=1060300 $Y=1096498
X4223 9037 8913 26 8973 25 8979 AOI21X1 $T=1070880 1089370 1 180 $X=1068580 $Y=1089118
X4224 9048 9100 26 8977 25 9236 AOI21X1 $T=1077320 1081990 1 0 $X=1077318 $Y=1078050
X4225 9130 9139 26 9114 25 9105 AOI21X1 $T=1079620 1059850 0 180 $X=1077320 $Y=1055910
X4226 9090 9132 26 9196 25 9080 AOI21X1 $T=1081000 1177930 0 0 $X=1080998 $Y=1177678
X4227 9097 9006 26 9197 25 9122 AOI21X1 $T=1081000 1229590 1 0 $X=1080998 $Y=1225650
X4228 9324 9248 26 9139 25 9140 AOI21X1 $T=1087900 1059850 1 180 $X=1085600 $Y=1059598
X4229 9254 9199 26 9290 25 9299 AOI21X1 $T=1087900 1089370 1 0 $X=1087898 $Y=1085430
X4230 9427 9373 26 9347 25 9220 AOI21X1 $T=1095720 1089370 0 180 $X=1093420 $Y=1085430
X4231 9277 9260 26 9377 25 9342 AOI21X1 $T=1093880 1185310 1 0 $X=1093878 $Y=1181370
X4232 9338 9248 26 9312 25 9474 AOI21X1 $T=1095720 1052470 0 0 $X=1095718 $Y=1052218
X4233 9520 9568 26 9530 25 9552 AOI21X1 $T=1105380 1045090 1 180 $X=1103080 $Y=1044838
X4234 9726 9707 26 9577 25 9677 AOI21X1 $T=1112280 1059850 0 180 $X=1109980 $Y=1055910
X4235 9829 9725 26 9568 25 9471 AOI21X1 $T=1113200 1045090 1 180 $X=1110900 $Y=1044838
X4236 9772 9862 26 9707 25 9819 AOI21X1 $T=1118260 1059850 1 0 $X=1118258 $Y=1055910
X4237 10016 9725 26 9869 25 9849 AOI21X1 $T=1121480 1037710 1 180 $X=1119180 $Y=1037458
X4238 9755 9899 26 9807 25 9850 AOI21X1 $T=1120560 1207450 1 0 $X=1120558 $Y=1203510
X4239 10201 10200 26 10179 25 9714 AOI21X1 $T=1135280 1037710 1 180 $X=1132980 $Y=1037458
X4240 10083 10189 26 10217 25 10140 AOI21X1 $T=1133900 1192690 1 0 $X=1133898 $Y=1188750
X4241 11454 11343 26 11438 25 11432 AOI21X1 $T=1200140 1332910 1 180 $X=1197840 $Y=1332658
X4242 181 11397 26 183 25 11580 AOI21X1 $T=1198300 1347670 0 0 $X=1198298 $Y=1347418
X4243 11741 11606 26 11754 25 205 AOI21X1 $T=1213480 1347670 1 0 $X=1213478 $Y=1343730
X4244 11848 11764 26 11776 25 11809 AOI21X1 $T=1217620 1096750 1 180 $X=1215320 $Y=1096498
X4245 12161 12209 26 12342 25 12377 AOI21X1 $T=1241080 1096750 1 0 $X=1241078 $Y=1092810
X4246 12449 12350 26 12329 25 12241 AOI21X1 $T=1243840 1052470 1 180 $X=1241540 $Y=1052218
X4247 12512 12381 26 12355 25 9250 AOI21X1 $T=1245220 1081990 0 180 $X=1242920 $Y=1078050
X4248 12347 12008 26 12547 25 12700 AOI21X1 $T=1249820 1170550 1 0 $X=1249818 $Y=1166610
X4249 12594 12650 26 12671 25 12535 AOI21X1 $T=1255340 1059850 0 0 $X=1255338 $Y=1059598
X4250 12849 12707 26 12717 25 12708 AOI21X1 $T=1260860 1104130 0 180 $X=1258560 $Y=1100190
X4251 12988 13003 26 13013 25 12552 AOI21X1 $T=1270980 1081990 1 0 $X=1270978 $Y=1078050
X4252 12582 13346 26 13386 25 13353 AOI21X1 $T=1288460 1155790 0 0 $X=1288458 $Y=1155538
X4253 13381 13236 26 13216 25 13486 AOI21X1 $T=1293520 1059850 0 0 $X=1293518 $Y=1059598
X4254 13451 13532 26 13553 25 10096 AOI21X1 $T=1297200 1067230 0 0 $X=1297198 $Y=1066978
X4255 13546 13588 26 13620 25 13477 AOI21X1 $T=1301340 1096750 1 0 $X=1301338 $Y=1092810
X4256 13631 13621 26 13597 25 13596 AOI21X1 $T=1304100 1118890 0 180 $X=1301800 $Y=1114950
X4257 9840 11527 26 11515 10484 25 11453 AOI22X1 $T=1203820 1185310 0 180 $X=1201060 $Y=1181370
X4258 9988 11849 26 11717 9920 25 11772 AOI22X1 $T=1218080 1163170 1 180 $X=1215320 $Y=1162918
X4259 9840 12268 26 12254 10484 25 12269 AOI22X1 $T=1239700 1155790 0 180 $X=1236940 $Y=1151850
X4260 9840 12563 26 12443 10484 25 12507 AOI22X1 $T=1252580 1133650 0 180 $X=1249820 $Y=1129710
X4261 9840 12779 26 12282 10484 25 12624 AOI22X1 $T=1262240 1126270 1 180 $X=1259480 $Y=1126018
X4262 9840 12794 26 12690 10484 25 12741 AOI22X1 $T=1262700 1111510 1 180 $X=1259940 $Y=1111258
X4263 9840 12919 26 12292 10484 25 12518 AOI22X1 $T=1269140 1111510 0 180 $X=1266380 $Y=1107570
X4264 9988 12873 26 12683 10484 25 13088 AOI22X1 $T=1267300 1052470 0 0 $X=1267298 $Y=1052218
X4265 9988 12940 26 12450 10484 25 12894 AOI22X1 $T=1270060 1074610 1 180 $X=1267300 $Y=1074358
X4266 9988 13022 26 12451 10484 25 12913 AOI22X1 $T=1273740 1096750 0 180 $X=1270980 $Y=1092810
X4267 9840 13036 26 12428 10484 25 13002 AOI22X1 $T=1274200 1067230 1 180 $X=1271440 $Y=1066978
X4268 9840 13121 26 11498 10484 25 13048 AOI22X1 $T=1278340 1081990 1 180 $X=1275580 $Y=1081738
X4269 9988 13122 26 12390 10484 25 13133 AOI22X1 $T=1276960 1096750 1 0 $X=1276958 $Y=1092810
X4270 9840 13163 26 12429 10484 25 13143 AOI22X1 $T=1279720 1081990 0 180 $X=1276960 $Y=1078050
X4271 9840 13164 26 12402 10484 25 13144 AOI22X1 $T=1279720 1089370 0 180 $X=1276960 $Y=1085430
X4272 9010 8874 25 8981 26 NAND2BX1 $T=1070880 1214830 0 180 $X=1069040 $Y=1210890
X4273 8911 8946 25 9078 26 NAND2BX1 $T=1069500 1163170 1 0 $X=1069498 $Y=1159230
X4274 9078 8920 25 9217 26 NAND2BX1 $T=1082380 1155790 1 0 $X=1082378 $Y=1151850
X4275 9217 8859 25 9264 26 NAND2BX1 $T=1086060 1148410 0 0 $X=1086058 $Y=1148158
X4276 9264 8677 25 9341 26 NAND2BX1 $T=1087900 1155790 1 0 $X=1087898 $Y=1151850
X4277 8736 9283 25 9108 26 NAND2BX1 $T=1089740 1222210 0 180 $X=1087900 $Y=1218270
X4278 9249 9241 25 9414 26 NAND2BX1 $T=1092960 1074610 1 0 $X=1092958 $Y=1070670
X4279 9341 8741 25 9282 26 NAND2BX1 $T=1093420 1155790 1 0 $X=1093418 $Y=1151850
X4280 9401 9501 25 9581 26 NAND2BX1 $T=1103540 1052470 1 0 $X=1103538 $Y=1048530
X4281 9596 9582 25 9883 26 NAND2BX1 $T=1112280 1067230 0 0 $X=1112278 $Y=1066978
X4282 9688 9621 25 9810 26 NAND2BX1 $T=1113200 1074610 1 0 $X=1113198 $Y=1070670
X4283 9784 9818 25 9887 26 NAND2BX1 $T=1122400 1059850 0 0 $X=1122398 $Y=1059598
X4284 9752 9835 25 10036 26 NAND2BX1 $T=1122860 1059850 1 0 $X=1122858 $Y=1055910
X4285 92 10047 25 10052 26 NAND2BX1 $T=1127460 1296010 0 0 $X=1127458 $Y=1295758
X4286 10073 10109 25 10218 26 NAND2BX1 $T=1129760 1200070 1 0 $X=1129758 $Y=1196130
X4287 10294 10276 25 10277 26 NAND2BX1 $T=1139880 1052470 1 180 $X=1138040 $Y=1052218
X4288 81 9915 74 25 26 9821 OA21XL $T=1123320 1303390 1 180 $X=1121020 $Y=1303138
X4289 10523 115 122 25 26 10670 OA21XL $T=1155520 1347670 0 0 $X=1155518 $Y=1347418
X4290 10523 10613 122 25 26 10729 OA21XL $T=1156440 1347670 1 0 $X=1156438 $Y=1343730
X4291 13326 13248 13298 25 26 12703 OA21XL $T=1287080 1170550 0 180 $X=1284780 $Y=1166610
X4292 34 39 9396 25 26 XNOR2XL $T=1094340 1347670 0 0 $X=1094338 $Y=1347418
X4293 28 53 9567 25 26 XNOR2XL $T=1102620 1347670 1 0 $X=1102618 $Y=1343730
X4294 9248 9391 9592 25 26 XNOR2XL $T=1103540 1059850 0 0 $X=1103538 $Y=1059598
X4295 28 83 86 25 26 XNOR2XL $T=1119640 1347670 0 0 $X=1119638 $Y=1347418
X4296 92 9871 9923 25 26 XNOR2XL $T=1124700 1296010 0 180 $X=1121480 $Y=1292070
X4297 9899 9901 9962 25 26 XNOR2XL $T=1121940 1200070 0 0 $X=1121938 $Y=1199818
X4298 34 90 93 25 26 XNOR2XL $T=1122860 1347670 0 0 $X=1122858 $Y=1347418
X4299 9862 10036 10093 25 26 XNOR2XL $T=1127920 1059850 1 0 $X=1127918 $Y=1055910
X4300 10189 10138 10094 25 26 XNOR2XL $T=1132060 1177930 0 180 $X=1128840 $Y=1173990
X4301 9725 10741 10762 25 26 XNOR2XL $T=1161960 1045090 0 0 $X=1161958 $Y=1044838
X4302 168 11305 11325 25 26 XNOR2XL $T=1190940 1332910 1 0 $X=1190938 $Y=1328970
X4303 11561 11546 11527 25 26 XNOR2XL $T=1205200 1185310 1 180 $X=1201980 $Y=1185058
X4304 12131 12149 11979 25 26 XNOR2XL $T=1233720 1118890 0 180 $X=1230500 $Y=1114950
X4305 13516 13500 12779 25 26 XNOR2XL $T=1297660 1126270 1 180 $X=1294440 $Y=1126018
X4306 9436 9375 25 9350 26 9328 NAND3BXL $T=1095720 1236970 1 180 $X=1093420 $Y=1236718
X4307 9438 9375 25 9417 26 9407 NAND3BXL $T=1098940 1236970 0 180 $X=1096640 $Y=1233030
X4308 9438 9417 25 9510 26 9814 NAND3BXL $T=1104460 1236970 0 0 $X=1104458 $Y=1236718
X4309 92 9382 25 9871 26 9851 NAND3BXL $T=1122860 1296010 1 180 $X=1120560 $Y=1295758
X4310 9871 92 25 9382 26 10292 NAND3BXL $T=1135740 1296010 0 0 $X=1135738 $Y=1295758
X4311 9107 9121 9128 26 25 9229 AOI2BB1X1 $T=1077320 1155790 0 0 $X=1077318 $Y=1155538
X4312 9636 9743 8947 26 25 9574 AOI2BB1X1 $T=1114120 1177930 0 180 $X=1111820 $Y=1173990
X4313 9636 9790 8827 26 25 9825 AOI2BB1X1 $T=1115040 1141030 1 0 $X=1115038 $Y=1137090
X4314 9740 10072 9243 26 25 9911 AOI2BB1X1 $T=1130220 1126270 1 180 $X=1127920 $Y=1126018
X4315 9740 10258 9437 26 25 10278 AOI2BB1X1 $T=1140340 1141030 0 180 $X=1138040 $Y=1137090
X4316 9740 10272 9518 26 25 10182 AOI2BB1X1 $T=1140340 1148410 1 180 $X=1138040 $Y=1148158
X4317 10417 10450 10435 26 25 10425 AOI2BB1X1 $T=1147240 1155790 1 180 $X=1144940 $Y=1155538
X4318 10417 10637 10602 26 25 10609 AOI2BB1X1 $T=1158280 1133650 1 180 $X=1155980 $Y=1133398
X4319 10417 11610 11425 26 25 11631 AOI2BB1X1 $T=1207040 1177930 1 0 $X=1207038 $Y=1173990
X4320 10417 11660 11561 26 25 11536 AOI2BB1X1 $T=1210720 1177930 1 180 $X=1208420 $Y=1177678
X4321 10417 11913 11314 26 25 11825 AOI2BB1X1 $T=1221760 1155790 1 180 $X=1219460 $Y=1155538
X4322 10417 11917 11449 26 25 11792 AOI2BB1X1 $T=1220840 1133650 0 0 $X=1220838 $Y=1133398
X4323 10417 12066 11345 26 25 12028 AOI2BB1X1 $T=1228660 1133650 0 180 $X=1226360 $Y=1129710
X4324 10417 12265 11220 26 25 12036 AOI2BB1X1 $T=1239700 1148410 0 180 $X=1237400 $Y=1144470
X4325 12364 12628 12622 26 25 12467 AOI2BB1X1 $T=1255800 1126270 0 180 $X=1253500 $Y=1122330
X4326 12364 12625 12514 26 25 12725 AOI2BB1X1 $T=1253960 1177930 1 0 $X=1253958 $Y=1173990
X4327 12364 12709 12463 26 25 12537 AOI2BB1X1 $T=1260860 1133650 1 180 $X=1258560 $Y=1133398
X4328 12364 12757 12744 26 25 12638 AOI2BB1X1 $T=1261320 1126270 0 180 $X=1259020 $Y=1122330
X4329 12364 12891 12874 26 25 12615 AOI2BB1X1 $T=1268220 1163170 0 180 $X=1265920 $Y=1159230
X4330 12364 12882 12889 26 25 12497 AOI2BB1X1 $T=1268680 1141030 1 180 $X=1266380 $Y=1140778
X4331 12364 12854 12926 26 25 12494 AOI2BB1X1 $T=1270060 1111510 1 180 $X=1267760 $Y=1111258
X4332 12364 12942 12927 26 25 12723 AOI2BB1X1 $T=1270060 1133650 1 180 $X=1267760 $Y=1133398
X4333 10046 10147 25 26 BUFX2 $T=1129300 1281250 0 0 $X=1129298 $Y=1280998
X4334 10495 10472 25 26 BUFX2 $T=1149540 1296010 0 0 $X=1149538 $Y=1295758
X4335 11728 11063 25 26 BUFX2 $T=1241540 1185310 1 0 $X=1241538 $Y=1181370
X4336 8875 25 8874 8875 8912 8969 26 OAI22XL $T=1060300 1214830 1 0 $X=1060298 $Y=1210890
X4337 8932 25 8936 8940 9041 9071 26 OAI22XL $T=1069960 1185310 1 0 $X=1069958 $Y=1181370
X4338 9109 25 9122 9109 9094 9123 26 OAI22XL $T=1078700 1222210 0 180 $X=1076400 $Y=1218270
X4339 8947 25 9096 9080 8948 9131 26 OAI22XL $T=1077780 1185310 0 0 $X=1077778 $Y=1185058
X4340 9174 25 9129 9174 9207 9201 26 OAI22XL $T=1081920 1200070 0 0 $X=1081918 $Y=1199818
X4341 9239 25 9178 9239 9195 9333 26 OAI22XL $T=1086060 1214830 1 0 $X=1086058 $Y=1210890
X4342 10380 25 11222 11230 10426 11290 26 OAI22XL $T=1186340 1236970 1 0 $X=1186338 $Y=1233030
X4343 11991 25 12001 12005 12024 11785 26 OAI22XL $T=1224980 1303390 0 0 $X=1224978 $Y=1303138
X4344 11988 25 12001 12016 12039 11811 26 OAI22XL $T=1225440 1244350 0 0 $X=1225438 $Y=1244098
X4345 12119 25 12001 12016 12143 11863 26 OAI22XL $T=1230960 1229590 0 0 $X=1230958 $Y=1229338
X4346 12323 25 12001 12016 12516 12212 26 OAI22XL $T=1248440 1214830 1 0 $X=1248438 $Y=1210890
X4347 12515 25 12345 12515 12564 12692 26 OAI22XL $T=1251200 1177930 0 0 $X=1251198 $Y=1177678
X4348 12001 25 12599 12589 12016 12194 26 OAI22XL $T=1253960 1244350 1 180 $X=1251660 $Y=1244098
X4349 13394 25 13353 13394 13385 13298 26 OAI22XL $T=1291680 1155790 0 180 $X=1289380 $Y=1151850
X4350 9393 8871 25 9013 26 9364 AND3XL $T=1096640 1177930 1 180 $X=1094340 $Y=1177678
X4351 9830 25 9822 26 74 9700 NAND3XL $T=1117800 1310770 0 180 $X=1115960 $Y=1306830
X4352 12322 25 12184 26 12345 12403 NAND3XL $T=1241540 1177930 0 0 $X=1241538 $Y=1177678
X4353 8873 8885 25 8827 8917 8875 26 8822 OAI32X1 $T=1060300 1207450 1 0 $X=1060298 $Y=1203510
X4354 9197 9097 25 9006 9151 9109 26 8948 OAI32X1 $T=1086520 1229590 1 0 $X=1086518 $Y=1225650
X4355 12192 12154 25 11220 12393 12564 26 11177 OAI32X1 $T=1249360 1170550 0 0 $X=1249358 $Y=1170298
X4356 13386 12582 25 13346 12685 13394 26 12889 OAI32X1 $T=1294440 1155790 0 0 $X=1294438 $Y=1155538
X4357 9218 9208 9201 25 9195 26 OAI2BB1X1 $T=1084220 1207450 1 180 $X=1081920 $Y=1207198
X4358 11273 168 11150 25 11343 26 OAI2BB1X1 $T=1189560 1340290 0 0 $X=1189558 $Y=1340038
X4359 8793 8742 8748 8824 25 26 8879 AO22XL $T=1054320 1118890 1 0 $X=1054318 $Y=1114950
X4360 8737 8742 8748 8793 25 26 8971 AO22XL $T=1060300 1126270 0 0 $X=1060298 $Y=1126018
X4361 8883 8916 8864 8871 25 26 8836 AO22XL $T=1063060 1185310 1 180 $X=1060300 $Y=1185058
X4362 8792 8814 8816 8935 25 26 8905 AO22XL $T=1066280 1111510 1 180 $X=1063520 $Y=1111258
X4363 8749 8734 8737 8961 25 26 9093 AO22XL $T=1069040 1126270 1 0 $X=1069038 $Y=1122330
X4364 8935 8742 8748 9013 25 26 9107 AO22XL $T=1075940 1155790 1 0 $X=1075938 $Y=1151850
X4365 9013 9270 9386 8952 25 26 9348 AO22XL $T=1097100 1118890 0 180 $X=1094340 $Y=1114950
X4366 9297 25 9208 26 9178 9326 NAND3X1 $T=1089740 1207450 1 180 $X=1087900 $Y=1207198
X4367 10739 25 10542 26 10724 10967 NAND3X1 $T=1162420 1281250 1 180 $X=1160580 $Y=1280998
X4368 8857 25 8746 8747 8744 8963 26 NAND4X1 $T=1048800 1126270 0 180 $X=1046500 $Y=1122330
X4369 8924 25 8933 8937 8930 8967 26 NAND4X1 $T=1063060 1155790 0 0 $X=1063058 $Y=1155538
X4370 8825 25 9256 9262 9276 9330 26 NAND4X1 $T=1086980 1133650 1 0 $X=1086978 $Y=1129710
X4371 9388 25 9331 9247 9349 9479 26 NAND4X1 $T=1095720 1163170 0 180 $X=1093420 $Y=1159230
X4372 9559 25 9350 9510 9503 9493 26 NAND4X1 $T=1103080 1244350 1 180 $X=1100780 $Y=1244098
X4373 9585 25 54 9567 9396 9652 26 NAND4X1 $T=1105840 1347670 1 180 $X=1103540 $Y=1347418
X4374 9909 25 9924 9929 9953 9535 26 NAND4X1 $T=1121940 1303390 1 0 $X=1121938 $Y=1299450
X4375 11429 25 11070 11446 11453 11175 26 NAND4X1 $T=1197840 1192690 1 0 $X=1197838 $Y=1188750
X4376 11748 25 11603 11730 11723 11718 26 NAND4X1 $T=1214400 1296010 1 180 $X=1212100 $Y=1295758
X4377 11670 25 11747 11751 11772 11868 26 NAND4X1 $T=1213480 1170550 1 0 $X=1213478 $Y=1166610
X4378 11897 25 11829 11602 11801 11957 26 NAND4X1 $T=1217620 1266490 1 180 $X=1215320 $Y=1266238
X4379 11982 25 11986 11987 11920 11983 26 NAND4X1 $T=1224520 1229590 1 0 $X=1224518 $Y=1225650
X4380 11994 25 12261 12277 12269 12330 26 NAND4X1 $T=1238320 1155790 0 0 $X=1238318 $Y=1155538
X4381 12343 25 12351 12356 12332 12004 26 NAND4X1 $T=1242460 1222210 0 0 $X=1242458 $Y=1221958
X4382 12133 25 12461 12495 12518 12389 26 NAND4X1 $T=1248440 1126270 0 0 $X=1248438 $Y=1126018
X4383 12276 25 12462 12496 12507 12232 26 NAND4X1 $T=1248440 1141030 1 0 $X=1248438 $Y=1137090
X4384 12100 25 12597 12614 12624 12420 26 NAND4X1 $T=1253040 1148410 1 0 $X=1253038 $Y=1144470
X4385 12659 25 12752 12764 12741 12781 26 NAND4X1 $T=1259940 1141030 1 0 $X=1259938 $Y=1137090
X4386 13001 25 12848 12879 12871 12860 26 NAND4X1 $T=1268220 1318150 1 180 $X=1265920 $Y=1317898
X4387 12724 25 12862 12890 12913 12896 26 NAND4X1 $T=1266380 1155790 1 0 $X=1266378 $Y=1151850
X4388 12875 25 12996 12999 12894 12930 26 NAND4X1 $T=1270520 1170550 0 0 $X=1270518 $Y=1170298
X4389 12699 25 13023 13031 13048 13008 26 NAND4X1 $T=1272360 1163170 1 0 $X=1272358 $Y=1159230
X4390 12751 25 13101 13109 13002 12993 26 NAND4X1 $T=1276040 1118890 1 0 $X=1276038 $Y=1114950
X4391 13096 25 12984 13021 13124 12994 26 NAND4X1 $T=1276040 1251730 0 0 $X=1276038 $Y=1251478
X4392 12595 25 13111 13116 13133 12911 26 NAND4X1 $T=1276500 1126270 0 0 $X=1276498 $Y=1126018
X4393 12586 25 13134 13117 13088 13102 26 NAND4X1 $T=1278800 1148410 0 180 $X=1276500 $Y=1144470
X4394 12605 25 13123 13127 13143 12945 26 NAND4X1 $T=1276960 1111510 0 0 $X=1276958 $Y=1111258
X4395 12850 25 13263 13271 13144 13237 26 NAND4X1 $T=1283860 1133650 0 0 $X=1283858 $Y=1133398
X4396 9506 9358 26 9521 9393 25 9695 AOI2BB2XL $T=1104460 1148410 1 0 $X=1104458 $Y=1144470
X4397 9553 9686 26 35 44 25 9902 AOI2BB2XL $T=1117800 1251730 0 0 $X=1117798 $Y=1251478
X4398 10003 9686 26 65 44 25 9908 AOI2BB2XL $T=1124240 1236970 0 180 $X=1121480 $Y=1233030
X4399 9802 9686 26 73 9963 25 10049 AOI2BB2XL $T=1123780 1236970 0 0 $X=1123778 $Y=1236718
X4400 10300 9686 26 101 9963 25 10270 AOI2BB2XL $T=1141260 1207450 0 180 $X=1138500 $Y=1203510
X4401 10408 10273 26 97 9963 25 10442 AOI2BB2XL $T=1144020 1192690 0 0 $X=1144018 $Y=1192438
X4402 10539 9686 26 108 9775 25 10403 AOI2BB2XL $T=1147700 1214830 1 180 $X=1144940 $Y=1214578
X4403 9974 9686 26 113 9963 25 10421 AOI2BB2XL $T=1148160 1236970 1 180 $X=1145400 $Y=1236718
X4404 10420 9686 26 94 9963 25 10540 AOI2BB2XL $T=1145860 1259110 0 0 $X=1145858 $Y=1258858
X4405 10703 10273 26 119 9963 25 10601 AOI2BB2XL $T=1160580 1200070 0 180 $X=1157820 $Y=1196130
X4406 10704 10273 26 127 9963 25 10937 AOI2BB2XL $T=1163800 1192690 0 0 $X=1163798 $Y=1192438
X4407 10969 10273 26 145 9775 25 10830 AOI2BB2XL $T=1174840 1296010 0 180 $X=1172080 $Y=1292070
X4408 10986 10273 26 132 9963 25 10949 AOI2BB2XL $T=1176220 1222210 0 180 $X=1173460 $Y=1218270
X4409 10122 10986 26 10067 149 25 10954 AOI2BB2XL $T=1176220 1236970 0 180 $X=1173460 $Y=1233030
X4410 10147 10987 26 10869 150 25 10955 AOI2BB2XL $T=1176220 1266490 0 180 $X=1173460 $Y=1262550
X4411 11025 10273 26 128 9963 25 10968 AOI2BB2XL $T=1177140 1266490 1 180 $X=1174380 $Y=1266238
X4412 10987 10273 26 130 9963 25 11130 AOI2BB2XL $T=1178980 1251730 1 0 $X=1178978 $Y=1247790
X4413 10122 11108 26 10067 160 25 11227 AOI2BB2XL $T=1179900 1214830 1 0 $X=1179898 $Y=1210890
X4414 11091 10273 26 133 9963 25 11095 AOI2BB2XL $T=1182660 1192690 1 180 $X=1179900 $Y=1192438
X4415 11108 10273 26 136 9963 25 11263 AOI2BB2XL $T=1180360 1214830 0 0 $X=1180358 $Y=1214578
X4416 11060 10273 26 155 9963 25 11148 AOI2BB2XL $T=1180360 1288630 1 0 $X=1180358 $Y=1284690
X4417 11188 10273 26 131 9963 25 11113 AOI2BB2XL $T=1183580 1244350 0 180 $X=1180820 $Y=1240410
X4418 11162 10273 26 135 9963 25 11110 AOI2BB2XL $T=1183580 1259110 0 180 $X=1180820 $Y=1255170
X4419 11228 10273 26 154 9504 25 11115 AOI2BB2XL $T=1183580 1296010 1 180 $X=1180820 $Y=1295758
X4420 10122 11188 26 10067 164 25 11251 AOI2BB2XL $T=1184040 1251730 1 0 $X=1184038 $Y=1247790
X4421 10122 11229 26 10067 163 25 11204 AOI2BB2XL $T=1188180 1222210 0 180 $X=1185420 $Y=1218270
X4422 11186 10273 26 175 9963 25 11161 AOI2BB2XL $T=1191860 1200070 1 180 $X=1189100 $Y=1199818
X4423 11324 10273 26 176 9775 25 11277 AOI2BB2XL $T=1192320 1296010 1 180 $X=1189560 $Y=1295758
X4424 11229 10273 26 157 9963 25 11381 AOI2BB2XL $T=1190940 1222210 1 0 $X=1190938 $Y=1218270
X4425 11335 10273 26 152 9963 25 11209 AOI2BB2XL $T=1193700 1229590 1 180 $X=1190940 $Y=1229338
X4426 11416 10273 26 123 9963 25 11307 AOI2BB2XL $T=1193700 1236970 0 180 $X=1190940 $Y=1233030
X4427 9652 10455 26 114 115 10428 25 NOR4BX1 $T=1146320 1347670 0 0 $X=1146318 $Y=1347418
X4428 8950 8941 8938 25 26 8924 AND3X2 $T=1065360 1133650 1 180 $X=1063060 $Y=1133398
X4429 12939 13026 13037 25 26 12932 AND3X2 $T=1272360 1318150 1 0 $X=1272358 $Y=1314210
X4430 8964 26 8931 8981 25 9007 9178 AOI211X1 $T=1075940 1207450 0 0 $X=1075938 $Y=1207198
X4431 9479 26 9393 9584 25 9599 9650 AOI211X1 $T=1104460 1155790 1 0 $X=1104458 $Y=1151850
X4432 9643 26 9665 9676 25 9435 9698 AOI211X1 $T=1109060 1214830 0 0 $X=1109058 $Y=1214578
X4433 9658 26 9393 9825 25 9838 9921 AOI211X1 $T=1116420 1133650 1 0 $X=1116418 $Y=1129710
X4434 8963 26 9393 9911 25 9764 9934 AOI211X1 $T=1121020 1126270 0 0 $X=1121018 $Y=1126018
X4435 8967 26 10176 10182 25 10118 10264 AOI211X1 $T=1132520 1155790 1 0 $X=1132518 $Y=1151850
X4436 9263 26 9393 10278 25 10180 10416 AOI211X1 $T=1137580 1133650 0 0 $X=1137578 $Y=1133398
X4437 9704 26 10176 10062 25 10283 10304 AOI211X1 $T=1138040 1177930 1 0 $X=1138038 $Y=1173990
X4438 9244 26 10176 10425 25 10303 10494 AOI211X1 $T=1144480 1163170 1 0 $X=1144478 $Y=1159230
X4439 9330 26 9393 10609 25 10604 10712 AOI211X1 $T=1155060 1133650 1 0 $X=1155058 $Y=1129710
X4440 10176 26 11445 11536 25 11548 11429 AOI211X1 $T=1202900 1177930 0 0 $X=1202898 $Y=1177678
X4441 10176 26 11585 11631 25 11526 11670 AOI211X1 $T=1207960 1170550 0 0 $X=1207958 $Y=1170298
X4442 10176 26 11617 11792 25 11545 11905 AOI211X1 $T=1214860 1141030 0 0 $X=1214858 $Y=1140778
X4443 10176 26 11750 11825 25 11726 11994 AOI211X1 $T=1215780 1148410 0 0 $X=1215778 $Y=1148158
X4444 10176 26 11945 12036 25 12022 12100 AOI211X1 $T=1225900 1148410 1 0 $X=1225898 $Y=1144470
X4445 10176 26 11560 12028 25 12065 12133 AOI211X1 $T=1226360 1126270 0 0 $X=1226358 $Y=1126018
X4446 10176 26 11589 12123 25 12092 12276 AOI211X1 $T=1231420 1141030 1 0 $X=1231418 $Y=1137090
X4447 10176 26 11777 12467 25 12499 12595 AOI211X1 $T=1247980 1126270 1 0 $X=1247978 $Y=1122330
X4448 10176 26 11778 12494 25 12517 12605 AOI211X1 $T=1248440 1111510 0 0 $X=1248438 $Y=1111258
X4449 10176 26 11413 12497 25 12064 12586 AOI211X1 $T=1248440 1141030 0 0 $X=1248438 $Y=1140778
X4450 10176 26 11902 12537 25 12132 12659 AOI211X1 $T=1249820 1133650 0 0 $X=1249818 $Y=1133398
X4451 10176 26 11618 12615 25 12583 12699 AOI211X1 $T=1253040 1163170 1 0 $X=1253038 $Y=1159230
X4452 10176 26 11722 12629 25 12639 12724 AOI211X1 $T=1253960 1155790 1 0 $X=1253958 $Y=1151850
X4453 10176 26 11727 12638 25 12648 12751 AOI211X1 $T=1254420 1118890 0 0 $X=1254418 $Y=1118638
X4454 10176 26 11861 12723 25 12674 12850 AOI211X1 $T=1258560 1133650 1 0 $X=1258558 $Y=1129710
X4455 10176 26 11643 12725 25 12621 12875 AOI211X1 $T=1258560 1170550 1 0 $X=1258558 $Y=1166610
X4456 9723 9687 25 9747 9547 9681 26 NAND4BX1 $T=1114580 1310770 1 180 $X=1111820 $Y=1310518
X4457 9880 9659 25 9896 9907 9372 26 NAND4BX1 $T=1120100 1192690 1 0 $X=1120098 $Y=1188750
X4458 9917 9921 25 9811 9951 9744 26 NAND4BX1 $T=1121940 1133650 0 0 $X=1121938 $Y=1133398
X4459 9889 9778 25 9910 9969 9801 26 NAND4BX1 $T=1122400 1111510 0 0 $X=1122398 $Y=1111258
X4460 10043 9679 25 10029 10064 9781 26 NAND4BX1 $T=1127460 1170550 1 0 $X=1127458 $Y=1166610
X4461 10034 9424 25 10038 10078 10107 26 NAND4BX1 $T=1127920 1118890 0 0 $X=1127918 $Y=1118638
X4462 10079 9650 25 9990 10066 9992 26 NAND4BX1 $T=1129300 1148410 0 0 $X=1129298 $Y=1148158
X4463 10150 9906 25 10119 10108 9966 26 NAND4BX1 $T=1132060 1141030 0 180 $X=1129300 $Y=1137090
X4464 10240 9799 25 10268 10282 10269 26 NAND4BX1 $T=1137120 1163170 0 0 $X=1137118 $Y=1162918
X4465 10259 9697 25 9885 10284 9967 26 NAND4BX1 $T=1137120 1185310 1 0 $X=1137118 $Y=1181370
X4466 10236 10304 25 10183 10325 10352 26 NAND4BX1 $T=1138960 1177930 0 0 $X=1138958 $Y=1177678
X4467 10527 9934 25 10434 10467 10448 26 NAND4BX1 $T=1149080 1133650 0 180 $X=1146320 $Y=1129710
X4468 10491 10416 25 10478 10468 10449 26 NAND4BX1 $T=1149080 1141030 0 180 $X=1146320 $Y=1137090
X4469 10614 10264 25 10625 10638 10532 26 NAND4BX1 $T=1155980 1155790 1 0 $X=1155978 $Y=1151850
X4470 10738 10494 25 10733 10771 10837 26 NAND4BX1 $T=1162420 1163170 1 0 $X=1162418 $Y=1159230
X4471 10802 10712 25 10822 10831 10533 26 NAND4BX1 $T=1165180 1133650 1 0 $X=1165178 $Y=1129710
X4472 11822 11905 25 11909 11927 11942 26 NAND4BX1 $T=1219920 1148410 1 0 $X=1219918 $Y=1144470
X4473 12530 12549 25 12526 12662 12686 26 NAND4BX1 $T=1254880 1310770 0 0 $X=1254878 $Y=1310518
X4474 13126 13136 25 13131 13103 12893 26 NAND4BX1 $T=1277420 1296010 1 0 $X=1277418 $Y=1292070
X4475 8953 8999 9009 9040 26 25 9263 OR4X1 $T=1069500 1141030 1 0 $X=1069498 $Y=1137090
X4476 9011 9071 9131 9146 26 25 9244 OR4X1 $T=1077320 1170550 0 0 $X=1077318 $Y=1170298
X4477 9348 9261 9200 9093 26 25 9146 OR4X1 $T=1088820 1126270 0 180 $X=1086060 $Y=1122330
X4478 11718 11957 11983 12004 26 25 12078 OR4X1 $T=1223600 1266490 0 0 $X=1223598 $Y=1266238
X4479 12994 12893 12860 12686 26 25 12190 OR4X1 $T=1268220 1296010 0 180 $X=1265460 $Y=1292070
X4480 11306 11068 11290 26 25 11344 OR3X2 $T=1190940 1185310 1 0 $X=1190938 $Y=1181370
X4481 11354 11332 11109 26 25 11087 OR3X2 $T=1193700 1259110 1 180 $X=1190940 $Y=1258858
X4482 9258 26 9243 9081 25 9265 9208 AOI211XL $T=1089740 1200070 1 180 $X=1087440 $Y=1199818
X4483 9915 26 81 9723 25 79 9830 AOI211XL $T=1120100 1318150 0 180 $X=1117800 $Y=1314210
X4484 10032 26 9930 9723 25 72 9909 AOI211XL $T=1124240 1310770 0 180 $X=1121940 $Y=1306830
X4485 9924 26 81 9930 25 88 9888 AOI211XL $T=1124240 1318150 1 180 $X=1121940 $Y=1317898
X4486 9363 9374 26 9376 9392 25 9402 9424 AOI221XL $T=1094340 1118890 0 0 $X=1094338 $Y=1118638
X4487 9573 9291 26 9734 9392 25 9684 9778 AOI221XL $T=1111820 1111510 1 0 $X=1111818 $Y=1107570
X4488 11744 188 26 11766 10448 25 11820 11782 AOI221XL $T=1213940 1214830 1 0 $X=1213938 $Y=1210890
X4489 11744 11504 26 11766 9801 25 11811 11831 AOI221XL $T=1213940 1244350 0 0 $X=1213938 $Y=1244098
X4490 11744 195 26 11766 10107 25 11841 11871 AOI221XL $T=1214860 1222210 0 0 $X=1214858 $Y=1221958
X4491 11744 203 26 11766 10352 25 11785 11773 AOI221XL $T=1218080 1310770 0 180 $X=1214860 $Y=1306830
X4492 11744 11562 26 11766 9992 25 11863 11783 AOI221XL $T=1215320 1229590 1 0 $X=1215318 $Y=1225650
X4493 11220 12154 26 11995 12183 25 12192 12322 AOI221XL $T=1232340 1177930 1 0 $X=1232338 $Y=1173990
X4494 11744 11246 26 10449 11766 25 12194 12220 AOI221XL $T=1232340 1244350 0 0 $X=1232338 $Y=1244098
X4495 11744 197 26 11766 10533 25 12212 12224 AOI221XL $T=1232800 1214830 1 0 $X=1232798 $Y=1210890
X4496 11744 245 26 11766 12330 25 12562 12505 AOI221XL $T=1254420 1340290 0 180 $X=1251200 $Y=1336350
X4497 11744 250 26 11766 11942 25 12607 12473 AOI221XL $T=1256260 1303390 0 180 $X=1253040 $Y=1299450
X4498 11744 257 26 11766 12420 25 12793 12819 AOI221XL $T=1259480 1340290 0 0 $X=1259478 $Y=1340038
X4499 11744 246 26 11766 12930 25 12944 12963 AOI221XL $T=1266840 1222210 0 0 $X=1266838 $Y=1221958
X4500 11744 244 26 11766 12945 25 12957 12985 AOI221XL $T=1267300 1273870 0 0 $X=1267298 $Y=1273618
X4501 11744 278 26 11766 12781 25 13046 13057 AOI221XL $T=1271440 1340290 1 0 $X=1271438 $Y=1336350
X4502 550 25 26 388 BUFX4 $T=1525360 1332910 1 0 $X=1525358 $Y=1328970
X4503 9419 44 41 25 26 9365 OAI2BB1XL $T=1096640 1332910 0 180 $X=1094340 $Y=1328970
X4504 28 44 43 25 26 9213 OAI2BB1XL $T=1096640 1347670 0 180 $X=1094340 $Y=1343730
X4505 9504 34 49 25 26 9087 OAI2BB1XL $T=1101700 1325530 1 180 $X=1099400 $Y=1325278
X4506 14400 14336 14377 13599 418 14270 14266 25 26 14214 14253 14235 13915 14214 14201 378 14123 3920 ICV_31 $T=1359300 1141030 1 180 $X=1350560 $Y=1140778
X4507 14465 14444 14568 13687 406 13744 14482 25 26 14475 14475 14445 365 14418 14394 398 14310 3920 ICV_31 $T=1375860 1229590 0 180 $X=1367120 $Y=1225650
X4508 14465 14482 14576 13687 417 14496 14488 25 26 14418 14436 14464 374 14239 14387 386 14245 3920 ICV_31 $T=1376780 1229590 1 180 $X=1368040 $Y=1229338
X4509 14150 14676 14577 396 438 14581 14549 25 26 14501 14561 14524 360 14489 14501 385 14484 3920 ICV_31 $T=1385520 1281250 1 180 $X=1376780 $Y=1280998
X4510 14400 14633 14748 13998 406 13906 14662 25 26 14661 14642 14571 14119 14595 14579 385 14547 3920 ICV_31 $T=1392420 1126270 0 180 $X=1383680 $Y=1122330
X4511 14465 14610 14765 13687 455 13660 14733 25 26 14715 14707 14686 381 14677 14632 386 14497 3920 ICV_31 $T=1400240 1251730 1 180 $X=1391500 $Y=1251478
X4512 14868 14770 14892 14865 469 14623 14816 25 26 14757 14807 14788 366 14758 14757 370 14435 3920 ICV_31 $T=1409900 1192690 0 180 $X=1401160 $Y=1188750
X4513 14751 14849 14836 14865 14596 14838 14817 25 26 14790 14812 14790 374 14745 14763 373 14328 3920 ICV_31 $T=1410360 1222210 1 180 $X=1401620 $Y=1221958
X4514 14607 14853 14932 14810 469 14671 14851 25 26 14789 14840 14818 354 14803 14789 13981 14229 3920 ICV_31 $T=1413120 1310770 0 180 $X=1404380 $Y=1306830
X4515 14607 14834 14970 14810 469 14581 14881 25 26 14793 14871 14813 361 14793 14780 377 14294 3920 ICV_31 $T=1417260 1281250 1 180 $X=1408520 $Y=1280998
X4516 15135 15289 15408 14865 15321 13875 15329 25 26 15327 15284 15288 371 15268 15252 373 15206 3920 ICV_31 $T=1461420 1222210 0 180 $X=1452680 $Y=1218270
X4517 15135 15371 15410 15340 515 13948 15331 25 26 15330 15218 15150 354 15170 15163 364 15207 3920 ICV_31 $T=1461880 1251730 0 180 $X=1453140 $Y=1247790
X4518 15292 15331 15414 15340 15321 13707 15335 25 26 15318 15330 15318 381 15280 15264 373 15223 3920 ICV_31 $T=1462340 1259110 1 180 $X=1453600 $Y=1258858
X4519 15353 15471 15454 14865 516 14731 15255 25 26 15322 15360 15327 371 15322 15287 373 15236 3920 ICV_31 $T=1468780 1214830 0 180 $X=1460040 $Y=1210890
X4520 15225 15477 15566 14810 515 14546 15489 25 26 15484 15484 15469 13853 15442 15433 523 15347 3920 ICV_31 $T=1479360 1325530 0 180 $X=1470620 $Y=1321590
X4521 15926 15872 15832 15687 511 14270 15777 25 26 15729 15770 15635 13879 15729 15714 401 15675 3920 ICV_31 $T=1507420 1133650 1 180 $X=1498680 $Y=1133398
X4522 15942 15897 15892 15340 515 14801 15827 25 26 15809 15756 15742 361 15732 15717 535 15726 3920 ICV_31 $T=1510640 1266490 0 180 $X=1501900 $Y=1262550
X4523 15926 15931 15930 15687 515 14663 15855 25 26 15850 15850 15836 13880 15799 15784 415 15571 3920 ICV_31 $T=1513860 1155790 0 180 $X=1505120 $Y=1151850
X4524 13560 13758 13768 11826 338 13374 13803 25 26 13894 13860 13877 13891 13557 13894 386 13968 3920 ICV_32 $T=1314680 1170550 0 0 $X=1314678 $Y=1170298
X4525 13640 13766 13773 13599 339 13734 13801 25 26 13868 13868 13659 13891 13852 13907 369 14025 3920 ICV_32 $T=1315140 1126270 0 0 $X=1315138 $Y=1126018
X4526 13609 13770 13777 11826 337 13712 13781 25 26 13896 13896 13887 366 13783 13903 378 13989 3920 ICV_32 $T=1315140 1192690 0 0 $X=1315138 $Y=1192438
X4527 13566 13771 13778 12746 338 13441 13733 25 26 13895 13844 13630 360 13655 13895 387 13984 3920 ICV_32 $T=1315140 1281250 0 0 $X=1315138 $Y=1280998
X4528 13081 13762 13776 12746 340 13741 13794 25 26 13888 13870 13888 13912 13765 13788 388 14000 3920 ICV_32 $T=1315140 1318150 0 0 $X=1315138 $Y=1317898
X4529 13560 13330 13787 13599 337 13735 13841 25 26 13897 13859 13460 13915 13317 13755 13883 14116 3920 ICV_32 $T=1315600 1163170 1 0 $X=1315598 $Y=1159230
X4530 348 349 13789 243 337 13890 13874 25 26 363 363 367 13853 380 383 378 13991 3920 ICV_32 $T=1315600 1347670 0 0 $X=1315598 $Y=1347418
X4531 13609 13781 13795 11826 338 13892 13822 25 26 13903 13896 13887 371 13783 13903 389 14011 3920 ICV_32 $T=1316060 1200070 1 0 $X=1316058 $Y=1196130
X4532 348 13747 13796 12746 340 13391 351 25 26 13889 13871 13889 13912 13368 13749 389 14015 3920 ICV_32 $T=1316980 1332910 0 0 $X=1316978 $Y=1332658
X4533 13349 13847 13823 13687 336 13746 13821 25 26 13929 13929 13637 361 13792 13963 389 14065 3920 ICV_32 $T=1320660 1244350 0 0 $X=1320658 $Y=1244098
X4534 13640 13855 13863 13599 342 13671 13766 25 26 13962 13753 13962 13915 14008 14001 364 14063 3920 ICV_32 $T=1322040 1141030 1 0 $X=1322038 $Y=1137090
X4535 13942 13951 13955 13599 342 13735 14094 25 26 14096 13897 13341 14119 13791 14137 385 14179 3920 ICV_32 $T=1331700 1163170 0 0 $X=1331698 $Y=1162918
X4536 13609 13952 13956 13998 338 13738 14088 25 26 14097 13997 13916 14119 13816 14097 378 14180 3920 ICV_32 $T=1331700 1207450 0 0 $X=1331698 $Y=1207198
X4537 13640 14024 14040 13599 342 13677 14047 25 26 14146 14147 14146 14119 14091 14208 385 14243 3920 ICV_32 $T=1337680 1118890 0 0 $X=1337678 $Y=1118638
X4538 12452 13985 13979 12746 362 13736 14002 25 26 14181 14173 14142 352 14181 14212 359 14258 3920 ICV_32 $T=1339980 1296010 1 0 $X=1339978 $Y=1292070
X4539 14599 14660 14666 396 455 13391 14683 25 26 14750 14750 14776 13893 14785 14798 13981 14309 3920 ICV_32 $T=1391500 1340290 1 0 $X=1391498 $Y=1336350
X4540 14599 15036 15044 14810 487 14546 15023 25 26 15137 15137 15157 13893 14934 15073 364 15250 3920 ICV_32 $T=1435660 1325530 1 0 $X=1435658 $Y=1321590
X4541 494 15041 15050 483 487 14391 15125 25 26 15134 15134 15151 13893 15166 15198 416 15271 3920 ICV_32 $T=1436120 1332910 0 0 $X=1436118 $Y=1332658
X4542 15358 15400 15404 14865 482 14586 15384 25 26 15505 15482 15505 13880 15235 15528 369 15564 3920 ICV_32 $T=1469240 1177930 1 0 $X=1469238 $Y=1173990
X4543 15135 15450 15451 15340 482 14405 15476 25 26 15576 15568 15576 374 15553 15597 536 15666 3920 ICV_32 $T=1478900 1244350 1 0 $X=1478898 $Y=1240410
X4544 13676 25 26 396 CLKINVX16 $T=1377700 1332910 0 0 $X=1377698 $Y=1332658
X4545 8885 26 8827 8873 25 8874 AOI21XL $T=1062600 1207450 1 180 $X=1060300 $Y=1207198
X4546 9127 26 9118 9092 25 9088 AOI21XL $T=1078700 1096750 0 180 $X=1076400 $Y=1092810
X4547 9534 26 9518 9502 25 9297 AOI21XL $T=1103080 1200070 0 180 $X=1100780 $Y=1196130
X4548 9477 26 9199 9373 25 9586 AOI21XL $T=1111820 1081990 0 0 $X=1111818 $Y=1081738
X4549 9904 26 9199 9927 25 9905 AOI21XL $T=1121480 1089370 1 0 $X=1121478 $Y=1085430
X4550 10228 26 9725 10200 25 10429 AOI21XL $T=1145400 1037710 0 0 $X=1145398 $Y=1037458
X4551 10732 26 9725 10865 25 10856 AOI21XL $T=1167020 1037710 0 0 $X=1167018 $Y=1037458
X4552 12231 26 12131 12157 25 12181 AOI21XL $T=1235560 1118890 1 180 $X=1233260 $Y=1118638
X4553 12152 26 12131 12209 25 12035 AOI21XL $T=1233720 1096750 0 0 $X=1233718 $Y=1096498
X4554 12588 26 12454 12672 25 12684 AOI21XL $T=1258560 1074610 0 180 $X=1256260 $Y=1070670
X4555 12253 26 11345 12630 25 12345 AOI21XL $T=1259480 1185310 0 0 $X=1259478 $Y=1185058
X4556 13586 26 13516 13613 25 13517 AOI21XL $T=1300880 1126270 0 0 $X=1300878 $Y=1126018
X4557 13651 26 13516 13621 25 13681 AOI21XL $T=1306400 1126270 0 0 $X=1306398 $Y=1126018
X4558 9426 45 25 26 INVX16 $T=1098940 1288630 1 180 $X=1094340 $Y=1288378
X4559 9746 70 25 26 INVX16 $T=1114580 1281250 1 180 $X=1109980 $Y=1280998
X4560 10418 111 25 26 INVX16 $T=1144020 1185310 1 0 $X=1144018 $Y=1181370
X4561 10443 100 25 26 INVX16 $T=1146780 1229590 1 0 $X=1146778 $Y=1225650
X4562 10857 109 25 26 INVX16 $T=1168400 1266490 0 0 $X=1168398 $Y=1266238
X4563 10799 139 25 26 INVX16 $T=1171620 1214830 0 0 $X=1171618 $Y=1214578
X4564 11090 143 25 26 INVX16 $T=1178980 1185310 1 0 $X=1178978 $Y=1181370
X4565 11821 227 25 26 INVX16 $T=1239240 1281250 1 0 $X=1239238 $Y=1277310
X4566 12259 231 25 26 INVX16 $T=1245680 1273870 0 180 $X=1241080 $Y=1269930
X4567 12458 213 25 26 INVX16 $T=1247520 1288630 1 0 $X=1247518 $Y=1284690
X4568 12548 235 25 26 INVX16 $T=1252580 1273870 0 180 $X=1247980 $Y=1269930
X4569 12405 242 25 26 INVX16 $T=1253040 1259110 0 180 $X=1248440 $Y=1255170
X4570 12221 241 25 26 INVX16 $T=1253500 1251730 1 180 $X=1248900 $Y=1251478
X4571 12596 264 25 26 INVX16 $T=1262240 1200070 0 0 $X=1262238 $Y=1199818
X4572 12876 280 25 26 INVX16 $T=1278340 1192690 0 0 $X=1278338 $Y=1192438
X4573 12877 279 25 26 INVX16 $T=1278340 1214830 1 0 $X=1278338 $Y=1210890
X4574 13233 289 25 26 INVX16 $T=1283860 1214830 1 180 $X=1279260 $Y=1214578
X4575 12780 284 25 26 INVX16 $T=1279720 1177930 0 0 $X=1279718 $Y=1177678
X4576 13227 300 25 26 INVX16 $T=1284780 1185310 0 0 $X=1284778 $Y=1185058
X4577 13293 321 25 26 INVX16 $T=1289380 1236970 0 0 $X=1289378 $Y=1236718
X4578 13387 309 25 26 INVX16 $T=1293060 1177930 0 0 $X=1293058 $Y=1177678
X4579 13563 308 25 26 INVX16 $T=1299960 1222210 1 0 $X=1299958 $Y=1218270
X4580 12134 11828 26 11437 12013 11147 25 11995 AOI32XL $T=1228200 1177930 0 180 $X=1224980 $Y=1173990
X4581 13174 13065 26 11344 13055 11243 25 13105 AOI32XL $T=1279720 1170550 1 180 $X=1276500 $Y=1170298
X4582 13325 12941 26 11225 12955 11087 25 13428 AOI32XL $T=1287540 1141030 0 0 $X=1287538 $Y=1140778
X4583 9108 9170 26 8732 9259 8736 25 9253 AOI32X1 $T=1085600 1214830 0 0 $X=1085598 $Y=1214578
X4584 9886 9952 26 9386 9918 9270 25 9748 AOI32X1 $T=1124240 1200070 0 180 $X=1121020 $Y=1196130
X4585 12703 12692 26 12403 12703 12753 25 9948 AOI32X1 $T=1258100 1177930 0 0 $X=1258098 $Y=1177678
X4586 13304 12815 26 11295 13010 11244 25 13247 AOI32X1 $T=1286620 1163170 1 180 $X=1283400 $Y=1162918
X4587 8883 9328 26 9354 9416 25 AOI2BB1XL $T=1092960 1229590 1 0 $X=1092958 $Y=1225650
X4588 9354 9522 26 8948 9676 25 AOI2BB1XL $T=1104460 1222210 1 0 $X=1104458 $Y=1218270
X4589 9636 9600 26 8870 9533 25 AOI2BB1XL $T=1106760 1163170 0 180 $X=1104460 $Y=1159230
X4590 9353 9358 26 9545 9569 25 AOI2BB1XL $T=1106760 1170550 1 180 $X=1104460 $Y=1170298
X4591 9636 9593 26 8940 9556 25 AOI2BB1XL $T=1106760 1192690 1 180 $X=1104460 $Y=1192438
X4592 9636 9716 26 8822 9736 25 AOI2BB1XL $T=1111360 1148410 1 0 $X=1111358 $Y=1144470
X4593 8871 9729 26 9740 9870 25 AOI2BB1XL $T=1111820 1192690 1 0 $X=1111818 $Y=1188750
X4594 9740 9839 26 8931 9769 25 AOI2BB1XL $T=1118720 1155790 1 180 $X=1116420 $Y=1155538
X4595 8748 9765 26 9740 9735 25 AOI2BB1XL $T=1119180 1133650 1 180 $X=1116880 $Y=1133398
X4596 9636 9895 26 8936 10062 25 AOI2BB1XL $T=1120560 1177930 1 0 $X=1120558 $Y=1173990
X4597 8961 9765 26 9740 9847 25 AOI2BB1XL $T=1122860 1118890 0 180 $X=1120560 $Y=1114950
X4598 8736 9729 26 9740 9754 25 AOI2BB1XL $T=1123320 1185310 0 180 $X=1121020 $Y=1181370
X4599 8749 9765 26 9740 9961 25 AOI2BB1XL $T=1121480 1155790 1 0 $X=1121478 $Y=1151850
X4600 8814 9729 26 9740 9912 25 AOI2BB1XL $T=1124240 1170550 1 180 $X=1121940 $Y=1170298
X4601 9930 9924 26 88 9822 25 AOI2BB1XL $T=1127000 1325530 1 0 $X=1126998 $Y=1321590
X4602 9003 9765 26 9740 9947 25 AOI2BB1XL $T=1129300 1126270 0 180 $X=1127000 $Y=1122330
X4603 8742 9729 26 9740 10137 25 AOI2BB1XL $T=1135740 1141030 1 180 $X=1133440 $Y=1140778
X4604 8816 9729 26 9740 10155 25 AOI2BB1XL $T=1135740 1170550 0 180 $X=1133440 $Y=1166610
X4605 8732 9991 26 9740 10101 25 AOI2BB1XL $T=1136200 1177930 1 180 $X=1133900 $Y=1177678
X4606 9101 9765 26 9740 10295 25 AOI2BB1XL $T=1141260 1126270 1 180 $X=1138960 $Y=1126018
X4607 9102 9765 26 10417 10565 25 AOI2BB1XL $T=1150000 1155790 1 0 $X=1149998 $Y=1151850
X4608 9228 9765 26 10417 10479 25 AOI2BB1XL $T=1153220 1148410 0 180 $X=1150920 $Y=1144470
X4609 9386 9729 26 10417 10647 25 AOI2BB1XL $T=1156440 1155790 0 0 $X=1156438 $Y=1155538
X4610 9270 9765 26 10417 10779 25 AOI2BB1XL $T=1163340 1141030 0 0 $X=1163338 $Y=1140778
X4611 11052 9729 26 10417 11590 25 AOI2BB1XL $T=1215320 1192690 0 180 $X=1213020 $Y=1188750
X4612 10967 9991 26 10417 11968 25 AOI2BB1XL $T=1225900 1155790 0 180 $X=1223600 $Y=1151850
X4613 11437 9729 26 10417 11914 25 AOI2BB1XL $T=1226360 1163170 1 180 $X=1224060 $Y=1162918
X4614 11147 9991 26 10417 12169 25 AOI2BB1XL $T=1231420 1155790 1 0 $X=1231418 $Y=1151850
X4615 10417 12153 26 11177 12123 25 AOI2BB1XL $T=1233720 1133650 1 180 $X=1231420 $Y=1133398
X4616 11322 9765 26 10417 12210 25 AOI2BB1XL $T=1232340 1126270 0 0 $X=1232338 $Y=1126018
X4617 11023 9991 26 12364 12438 25 AOI2BB1XL $T=1242920 1155790 1 0 $X=1242918 $Y=1151850
X4618 11323 9729 26 12364 12334 25 AOI2BB1XL $T=1245220 1141030 1 180 $X=1242920 $Y=1140778
X4619 11295 9765 26 12364 12623 25 AOI2BB1XL $T=1249820 1155790 0 0 $X=1249818 $Y=1155538
X4620 11344 9991 26 12364 12956 25 AOI2BB1XL $T=1258560 1163170 0 0 $X=1258558 $Y=1162918
X4621 12364 12710 26 12729 12629 25 AOI2BB1XL $T=1260860 1155790 1 180 $X=1258560 $Y=1155538
X4622 11275 9991 26 12364 12719 25 AOI2BB1XL $T=1259940 1155790 1 0 $X=1259938 $Y=1151850
X4623 11063 9729 26 12364 12920 25 AOI2BB1XL $T=1266840 1177930 0 0 $X=1266838 $Y=1177678
X4624 11066 9729 26 12364 13112 25 AOI2BB1XL $T=1279720 1155790 1 180 $X=1277420 $Y=1155538
X4625 11087 9729 26 12364 13059 25 AOI2BB1XL $T=1280180 1118890 1 180 $X=1277880 $Y=1118638
X4626 11225 9729 26 12364 13262 25 AOI2BB1XL $T=1282940 1126270 1 0 $X=1282938 $Y=1122330
X4627 11243 9729 26 12364 13241 25 AOI2BB1XL $T=1285240 1141030 1 180 $X=1282940 $Y=1140778
X4628 11244 9729 26 12364 13148 25 AOI2BB1XL $T=1285700 1126270 1 180 $X=1283400 $Y=1126018
X4629 10045 9994 25 9554 10125 26 10148 9097 OAI221X1 $T=1128840 1281250 1 0 $X=1128838 $Y=1277310
X4630 10045 10248 25 9782 10125 26 10307 9283 OAI221X1 $T=1137120 1273870 1 0 $X=1137118 $Y=1269930
X4631 10045 10296 25 10300 10125 26 10333 9238 OAI221X1 $T=1138040 1214830 1 0 $X=1138038 $Y=1210890
X4632 10045 9922 25 9418 10125 26 10444 9151 OAI221X1 $T=1143560 1273870 0 0 $X=1143558 $Y=1273618
X4633 10362 10546 25 10534 10125 26 10572 9509 OAI221X1 $T=1150000 1281250 1 0 $X=1149998 $Y=1277310
X4634 10045 11085 25 11091 10751 26 11121 10136 OAI221X1 $T=1178520 1200070 1 0 $X=1178518 $Y=1196130
X4635 10380 11289 25 11310 10426 26 11227 11421 OAI221X1 $T=1201060 1214830 0 180 $X=1197380 $Y=1210890
X4636 10888 10362 25 10669 10751 26 11911 11546 OAI221X1 $T=1218080 1281250 0 0 $X=1218078 $Y=1280998
X4637 10362 11111 25 11060 10751 26 12185 11926 OAI221X1 $T=1231420 1288630 1 0 $X=1231418 $Y=1284690
X4638 10362 11431 25 11324 10751 26 12189 11941 OAI221X1 $T=1231880 1288630 0 0 $X=1231878 $Y=1288378
X4639 10792 10362 25 10777 10751 26 12357 11901 OAI221X1 $T=1240620 1288630 0 0 $X=1240618 $Y=1288378
X4640 10362 11202 25 11162 10751 26 12587 12500 OAI221X1 $T=1249820 1251730 1 0 $X=1249818 $Y=1247790
X4641 10362 11336 25 10987 10751 26 12765 12857 OAI221X1 $T=1258100 1251730 0 0 $X=1258098 $Y=1251478
X4642 10362 11285 25 11416 10751 26 12777 12834 OAI221X1 $T=1258560 1236970 0 0 $X=1258558 $Y=1236718
X4643 10362 11374 25 11188 10751 26 12745 12730 OAI221X1 $T=1263160 1244350 1 180 $X=1259480 $Y=1244098
X4644 10362 11230 25 11335 10751 26 12816 12814 OAI221X1 $T=1259940 1229590 0 0 $X=1259938 $Y=1229338
X4645 10362 11310 25 11108 10751 26 12884 12929 OAI221X1 $T=1265000 1207450 0 0 $X=1264998 $Y=1207198
X4646 10362 11266 25 11186 10751 26 12937 12943 OAI221X1 $T=1266380 1207450 1 0 $X=1266378 $Y=1203510
X4647 8883 9151 25 26 9091 OR2XL $T=1080540 1236970 0 180 $X=1078700 $Y=1233030
X4648 8871 9097 25 26 9194 OR2XL $T=1086060 1192690 1 180 $X=1084220 $Y=1192438
X4649 9006 9097 25 26 9755 OR2XL $T=1112280 1207450 0 0 $X=1112278 $Y=1207198
X4650 9225 9509 25 26 10083 OR2XL $T=1127920 1192690 1 0 $X=1127918 $Y=1188750
X4651 10445 10166 25 26 10542 OR2XL $T=1146320 1288630 1 0 $X=1146318 $Y=1284690
X4652 10777 10147 25 26 10724 OR2XL $T=1163800 1288630 0 180 $X=1161960 $Y=1284690
X4653 11052 11546 25 26 11588 OR2XL $T=1205200 1118890 0 0 $X=1205198 $Y=1118638
X4654 11736 12641 25 26 12939 OR2XL $T=1260860 1310770 0 0 $X=1260858 $Y=1310518
X4655 10050 10045 25 9553 10125 10146 8885 26 OAI221X2 $T=1127460 1259110 1 0 $X=1127458 $Y=1255170
X4656 10074 10045 25 9802 10125 10165 9061 26 OAI221X2 $T=1128380 1236970 0 0 $X=1128378 $Y=1236718
X4657 10095 10045 25 10003 10125 10174 9138 26 OAI221X2 $T=1128840 1229590 1 0 $X=1128838 $Y=1225650
X4658 10265 10045 25 9699 10125 10334 8917 26 OAI221X2 $T=1136660 1266490 1 0 $X=1136658 $Y=1262550
X4659 10402 10045 25 10408 10125 10462 9258 26 OAI221X2 $T=1143100 1207450 0 0 $X=1143098 $Y=1207198
X4660 10571 10045 25 10539 10125 10611 9512 26 OAI221X2 $T=1151840 1222210 0 0 $X=1151838 $Y=1221958
X4661 10588 10045 25 10420 10125 10627 8964 26 OAI221X2 $T=1152760 1259110 1 0 $X=1152758 $Y=1255170
X4662 10454 10045 25 9974 10125 10635 8834 26 OAI221X2 $T=1153220 1236970 0 0 $X=1153218 $Y=1236718
X4663 10766 10045 25 10704 10751 10838 9806 26 OAI221X2 $T=1162880 1200070 1 0 $X=1162878 $Y=1196130
X4664 10626 10045 25 10703 10751 10839 9534 26 OAI221X2 $T=1162880 1200070 0 0 $X=1162878 $Y=1199818
X4665 10445 9929 25 10969 10147 10998 11023 26 OAI221X2 $T=1171620 1288630 1 0 $X=1171618 $Y=1284690
X4666 11114 10362 25 11025 10751 12283 12253 26 OAI221X2 $T=1235560 1266490 1 0 $X=1235558 $Y=1262550
X4667 11465 10362 25 11229 10751 12579 12582 26 OAI221X2 $T=1247980 1222210 1 0 $X=1247978 $Y=1218270
X4668 11216 10362 25 11228 10751 12661 12393 26 OAI221X2 $T=1252120 1288630 0 0 $X=1252118 $Y=1288378
X4669 10919 10362 25 10986 10751 12675 12685 26 OAI221X2 $T=1262240 1229590 0 180 $X=1257180 $Y=1225650
X4670 10791 10362 25 10969 10751 12711 12154 26 OAI221X2 $T=1263620 1288630 1 180 $X=1258560 $Y=1288378
X4671 9007 8964 25 8931 8834 8912 26 8870 OAI32XL $T=1068580 1200070 1 180 $X=1065360 $Y=1199818
X4672 8982 9138 25 9005 9061 9174 26 8880 OAI32XL $T=1078240 1207450 1 0 $X=1078238 $Y=1203510
X4673 9265 9258 25 9243 9238 9207 26 8980 OAI32XL $T=1088360 1200070 0 180 $X=1085140 $Y=1196130
X4674 9502 9534 25 9518 9512 9406 26 9437 OAI32XL $T=1102620 1200070 0 0 $X=1102618 $Y=1199818
X4675 12630 12253 25 11345 12500 12515 26 12463 OAI32XL $T=1251660 1185310 0 180 $X=1248440 $Y=1181370
X4676 10322 10490 10634 9916 10423 25 26 10742 MX3XL $T=1154600 1111510 1 0 $X=1154598 $Y=1107570
X4677 10331 10493 10787 9916 10397 25 26 10847 MX3XL $T=1161960 1096750 0 0 $X=1161958 $Y=1096498
X4678 10331 10615 10788 9916 10653 25 26 10848 MX3XL $T=1161960 1104130 1 0 $X=1161958 $Y=1100190
X4679 10207 10794 10930 10331 10465 25 26 10866 MX3XL $T=1175760 1111510 0 180 $X=1169780 $Y=1107570
X4680 10331 10787 10939 10887 10728 25 26 11057 MX3XL $T=1170240 1096750 0 0 $X=1170238 $Y=1096498
X4681 10716 10803 10892 140 10995 25 26 11005 MX3XL $T=1170700 1177930 1 0 $X=1170698 $Y=1173990
X4682 10207 10952 10945 10331 10536 25 26 10904 MX3XL $T=1176680 1096750 0 180 $X=1170700 $Y=1092810
X4683 10207 11007 10962 10322 10782 25 26 10921 MX3XL $T=1177600 1118890 1 180 $X=1171620 $Y=1118638
X4684 10951 10965 11004 11030 11056 25 26 11127 MX3XL $T=1173460 1045090 0 0 $X=1173458 $Y=1044838
X4685 10331 10788 11079 10887 11128 25 26 11144 MX3XL $T=1176680 1104130 1 0 $X=1176678 $Y=1100190
X4686 10951 11039 10928 11030 11153 25 26 11182 MX3XL $T=1178060 1067230 0 0 $X=1178058 $Y=1066978
X4687 11206 11190 11127 11133 11101 25 26 10323 MX3XL $T=1185880 1052470 0 180 $X=1179900 $Y=1048530
X4688 10207 10891 11143 10331 10551 25 26 11093 MX3XL $T=1185880 1089370 1 180 $X=1179900 $Y=1089118
X4689 10207 10962 11145 10322 10810 25 26 11094 MX3XL $T=1185880 1118890 1 180 $X=1179900 $Y=1118638
X4690 10951 11004 11160 11030 11205 25 26 11234 MX3XL $T=1180820 1037710 1 0 $X=1180818 $Y=1033770
X4691 10299 11219 11184 10207 10930 25 26 11062 MX3XL $T=1187720 1111510 1 180 $X=1181740 $Y=1111258
X4692 11030 11194 11082 11241 11265 25 26 11272 MX3XL $T=1184040 1074610 1 0 $X=1184038 $Y=1070670
X4693 11241 11274 11182 11133 11200 25 26 10186 MX3XL $T=1190940 1067230 1 180 $X=1184960 $Y=1066978
X4694 11030 11138 11194 11241 11330 25 26 11313 MX3XL $T=1187260 1067230 1 0 $X=1187258 $Y=1063290
X4695 10299 11320 11279 10207 11235 25 26 10939 MX3XL $T=1193240 1096750 1 180 $X=1187260 $Y=1096498
X4696 10299 11279 11280 10207 11236 25 26 11079 MX3XL $T=1193240 1104130 1 180 $X=1187260 $Y=1103878
X4697 11030 11142 10927 11206 11342 25 26 11350 MX3XL $T=1187720 1045090 0 0 $X=1187718 $Y=1044838
X4698 11030 10938 11038 11206 11250 25 26 11061 MX3XL $T=1193700 1037710 1 180 $X=1187720 $Y=1037458
X4699 10470 11425 11449 10299 11184 25 26 11145 MX3XL $T=1202440 1118890 1 180 $X=1196460 $Y=1118638
X4700 11030 11119 10994 11241 11534 25 26 11535 MX3XL $T=1198760 1059850 1 0 $X=1198758 $Y=1055910
X4701 11206 11565 11278 11133 11488 25 26 10065 MX3XL $T=1206580 1037710 0 180 $X=1200600 $Y=1033770
X4702 11241 11607 11190 11133 11529 25 26 10123 MX3XL $T=1208880 1052470 1 180 $X=1202900 $Y=1052218
X4703 11241 11912 11274 11242 11860 25 26 10550 MX3XL $T=1223140 1067230 0 180 $X=1217160 $Y=1063290
X4704 10536 10331 10548 10371 25 26 9916 10643 MXI3X1 $T=1150460 1096750 0 0 $X=1150458 $Y=1096498
X4705 10551 10331 10447 9777 25 26 9916 10706 MXI3X1 $T=1151380 1089370 0 0 $X=1151378 $Y=1089118
X4706 10810 10322 10624 10181 25 26 10887 10958 MXI3X1 $T=1165640 1118890 1 0 $X=1165638 $Y=1114950
X4707 8871 10470 8736 10928 25 26 10619 11082 MXI3X1 $T=1172540 1074610 0 0 $X=1172538 $Y=1074358
X4708 11062 10322 11051 10388 25 26 10887 11237 MXI3X1 $T=1178520 1118890 1 0 $X=1178518 $Y=1114950
X4709 11220 10764 11177 10870 25 26 10871 11083 MXI3X1 $T=1186800 1155790 0 180 $X=1179440 $Y=1151850
X4710 11213 10908 11088 11269 25 26 140 11346 MXI3X1 $T=1185880 1148410 1 0 $X=1185878 $Y=1144470
X4711 11425 10764 11314 11054 25 26 141 11223 MXI3X1 $T=1194160 1170550 0 180 $X=1186800 $Y=1166610
X4712 11177 10750 11345 11102 25 26 10871 11253 MXI3X1 $T=1195540 1133650 1 180 $X=1188180 $Y=1133398
X4713 11314 10764 11220 11031 25 26 10871 11213 MXI3X1 $T=1196460 1148410 1 180 $X=1189100 $Y=1148158
X4714 11265 11241 11398 11383 25 26 11133 9949 MXI3X1 $T=1198760 1074610 1 180 $X=1191400 $Y=1074358
X4715 11405 10716 11203 11321 25 26 140 11541 MXI3X1 $T=1196920 1148410 1 0 $X=1196918 $Y=1144470
X4716 11223 10716 11450 11198 25 26 140 11467 MXI3X1 $T=1196920 1170550 0 0 $X=1196918 $Y=1170298
X4717 11534 11241 11505 11485 25 26 11133 10754 MXI3X1 $T=1204280 1067230 1 180 $X=1196920 $Y=1066978
X4718 11330 11241 11608 11587 25 26 11133 10636 MXI3X1 $T=1210260 1074610 1 180 $X=1202900 $Y=1074358
X4719 11342 11241 11712 11690 25 26 11242 10966 MXI3X1 $T=1214400 1052470 0 180 $X=1207040 $Y=1048530
X4720 11250 11241 11867 11846 25 26 11242 10544 MXI3X1 $T=1220840 1045090 0 180 $X=1213480 $Y=1041150
X4721 10464 10266 10407 10263 25 26 MXI2XL $T=1148160 1089370 1 180 $X=1144940 $Y=1089118
X4722 8961 126 10756 9003 25 26 MXI2XL $T=1161040 1133650 1 0 $X=1161038 $Y=1129710
X4723 9270 126 10772 9386 25 26 MXI2XL $T=1161500 1170550 0 0 $X=1161498 $Y=1170298
X4724 8814 126 10776 8816 25 26 MXI2XL $T=1162420 1170550 1 0 $X=1162418 $Y=1166610
X4725 8742 10764 10753 8748 25 26 MXI2XL $T=1165640 1163170 1 180 $X=1162420 $Y=1162918
X4726 9003 10764 10811 9101 25 26 MXI2XL $T=1163340 1155790 0 0 $X=1163338 $Y=1155538
X4727 8736 10470 10832 8732 25 26 MXI2XL $T=1164260 1155790 1 0 $X=1164258 $Y=1151850
X4728 8749 10764 10853 8961 25 26 MXI2XL $T=1165180 1177930 1 0 $X=1165178 $Y=1173990
X4729 9101 126 10901 9228 25 26 MXI2XL $T=1167940 1141030 1 0 $X=1167938 $Y=1137090
X4730 8732 126 10947 8742 25 26 MXI2XL $T=1171620 1141030 0 0 $X=1171618 $Y=1140778
X4731 8748 126 10931 8814 25 26 MXI2XL $T=1174840 1148410 1 180 $X=1171620 $Y=1148158
X4732 8871 126 10963 8736 25 26 MXI2XL $T=1172540 1133650 0 0 $X=1172538 $Y=1133398
X4733 8816 126 10946 8749 25 26 MXI2XL $T=1175760 1126270 1 180 $X=1172540 $Y=1126018
X4734 9228 10764 10984 9102 25 26 MXI2XL $T=1173000 1163170 1 0 $X=1172998 $Y=1159230
X4735 9102 126 11067 9270 25 26 MXI2XL $T=1177140 1148410 0 0 $X=1177138 $Y=1148158
X4736 11063 10750 11102 11087 25 26 MXI2XL $T=1178060 1126270 0 0 $X=1178058 $Y=1126018
X4737 11066 10764 11125 11063 25 26 MXI2XL $T=1178980 1177930 1 0 $X=1178978 $Y=1173990
X4738 8883 10764 11120 8871 25 26 MXI2XL $T=1183580 1177930 1 180 $X=1180360 $Y=1177678
X4739 11173 140 11146 11076 25 26 MXI2XL $T=1184960 1170550 0 180 $X=1181740 $Y=1166610
X4740 9386 10470 11176 11066 25 26 MXI2XL $T=1184960 1126270 1 0 $X=1184958 $Y=1122330
X4741 11244 10764 11054 11295 25 26 MXI2XL $T=1187720 1163170 1 0 $X=1187718 $Y=1159230
X4742 11275 10764 11303 11322 25 26 MXI2XL $T=1189100 1177930 0 0 $X=1189098 $Y=1177678
X4743 11087 10764 10870 11225 25 26 MXI2XL $T=1192320 1155790 1 180 $X=1189100 $Y=1155538
X4744 11023 10470 11184 11147 25 26 MXI2XL $T=1190020 1118890 0 0 $X=1190018 $Y=1118638
X4745 11225 10764 11031 11244 25 26 MXI2XL $T=1193240 1155790 0 180 $X=1190020 $Y=1151850
X4746 11344 10750 11212 11275 25 26 MXI2XL $T=1193700 1126270 0 180 $X=1190480 $Y=1122330
X4747 11295 10764 11107 11243 25 26 MXI2XL $T=1196460 1155790 1 0 $X=1196458 $Y=1151850
X4748 11243 10764 10878 11344 25 26 MXI2XL $T=1199680 1177930 1 180 $X=1196460 $Y=1177678
X4749 11142 11389 11190 11506 25 26 MXI2XL $T=1196920 1045090 0 0 $X=1196918 $Y=1044838
X4750 11322 10470 11219 11323 25 26 MXI2XL $T=1201520 1118890 0 180 $X=1198300 $Y=1114950
X4751 8883 11242 11530 11483 25 26 MXI2XL $T=1201060 1126270 0 0 $X=1201058 $Y=1126018
X4752 11119 11389 11274 11613 25 26 MXI2XL $T=1205200 1059850 1 0 $X=1205198 $Y=1055910
X4753 9398 40 26 25 BUFX16 $T=1098020 1288630 0 180 $X=1091580 $Y=1284690
X4754 9526 51 26 25 BUFX16 $T=1103540 1251730 1 180 $X=1097100 $Y=1251478
X4755 9662 55 26 25 BUFX16 $T=1109980 1251730 0 180 $X=1103540 $Y=1247790
X4756 9767 56 26 25 BUFX16 $T=1117340 1266490 1 180 $X=1110900 $Y=1266238
X4757 10020 87 26 25 BUFX16 $T=1125160 1222210 1 180 $X=1118720 $Y=1221958
X4758 9996 80 26 25 BUFX16 $T=1125620 1214830 1 180 $X=1119180 $Y=1214578
X4759 10229 75 26 25 BUFX16 $T=1136660 1229590 1 180 $X=1130220 $Y=1229338
X4760 10645 117 26 25 BUFX16 $T=1157360 1229590 1 0 $X=1157358 $Y=1225650
X4761 10713 124 26 25 BUFX16 $T=1161040 1185310 1 0 $X=1161038 $Y=1181370
X4762 11364 177 26 25 BUFX16 $T=1204740 1281250 1 0 $X=1204738 $Y=1277310
X4763 10465 10322 10407 10120 25 26 9916 10594 MXI3XL $T=1147240 1111510 1 0 $X=1147238 $Y=1107570
X4764 10782 10322 10545 10400 25 26 10887 10917 MXI3XL $T=1164260 1118890 0 0 $X=1164258 $Y=1118638
X4765 10877 140 10918 8883 25 26 10908 11089 MXI3XL $T=1168860 1163170 0 0 $X=1168858 $Y=1162918
X4766 11052 126 10967 10948 25 26 141 10892 MXI3XL $T=1177140 1185310 0 180 $X=1169780 $Y=1181370
X4767 11135 173 11260 8951 25 26 10716 11413 MXI3XL $T=1189100 1141030 0 0 $X=1189098 $Y=1140778
X4768 11449 10764 11425 11107 25 26 10469 11405 MXI3XL $T=1204740 1148410 1 180 $X=1197380 $Y=1148158
X4769 9953 10445 11060 10147 11092 11147 25 26 OAI221X4 $T=1177600 1273870 0 0 $X=1177598 $Y=1273618
X4770 10380 10933 10919 10426 10954 11066 25 26 OAI221X4 $T=1178980 1236970 1 0 $X=1178978 $Y=1233030
X4771 10530 10445 11186 10122 11208 11243 25 26 OAI221X4 $T=1183580 1185310 0 0 $X=1183578 $Y=1185058
X4772 10595 10445 11162 10122 11238 11275 25 26 OAI221X4 $T=1185420 1200070 1 0 $X=1185418 $Y=1196130
X4773 10486 10445 11025 10122 11155 11322 25 26 OAI221X4 $T=1187720 1192690 0 0 $X=1187718 $Y=1192438
X4774 10924 10445 11228 10147 11276 11323 25 26 OAI221X4 $T=1187720 1281250 0 0 $X=1187718 $Y=1280998
X4775 10380 11289 11310 10426 11227 11244 25 26 OAI221X4 $T=1192780 1214830 0 180 $X=1187720 $Y=1210890
X4776 10380 11318 11374 10290 11251 11225 25 26 OAI221X4 $T=1195540 1251730 0 180 $X=1190480 $Y=1247790
X4777 9915 10445 11324 10147 11390 11437 25 26 OAI221X4 $T=1196000 1288630 0 0 $X=1195998 $Y=1288378
X4778 11406 10445 11416 10122 11353 11295 25 26 OAI221X4 $T=1196920 1192690 0 0 $X=1196918 $Y=1192438
X4779 8946 8940 8920 8936 25 26 9000 OA22XL $T=1068120 1163170 0 0 $X=1068118 $Y=1162918
X4780 8936 8943 9177 8822 25 26 9247 OA22XL $T=1081460 1163170 0 0 $X=1081458 $Y=1162918
X4781 8947 8677 8741 8940 25 26 9349 OA22XL $T=1085600 1155790 0 0 $X=1085598 $Y=1155538
X4782 8827 9141 9119 8870 25 26 9331 OA22XL $T=1087440 1163170 0 0 $X=1087438 $Y=1162918
X4783 8931 9353 9359 8880 25 26 9388 OA22XL $T=1093420 1163170 0 0 $X=1093418 $Y=1162918
X4784 10792 10290 10260 10743 25 26 10739 OA22XL $T=1166100 1288630 1 180 $X=1163340 $Y=1288378
X4785 10777 10273 85 10372 25 26 10735 OA22XL $T=1166100 1296010 0 180 $X=1163340 $Y=1292070
X4786 10290 11114 11103 10260 25 26 11155 OA22XL $T=1180360 1273870 1 0 $X=1180358 $Y=1269930
X4787 10290 11111 11122 10260 25 26 11092 OA22XL $T=1184040 1281250 0 180 $X=1181280 $Y=1277310
X4788 10290 11202 11163 10260 25 26 11238 OA22XL $T=1184960 1266490 1 0 $X=1184958 $Y=1262550
X4789 10426 11266 11187 10260 25 26 11208 OA22XL $T=1191400 1229590 0 180 $X=1188640 $Y=1225650
X4790 10426 11285 11291 10260 25 26 11353 OA22XL $T=1189560 1244350 1 0 $X=1189558 $Y=1240410
X4791 10290 11216 11210 10260 25 26 11276 OA22XL $T=1192320 1288630 1 180 $X=1189560 $Y=1288378
X4792 11316 11206 11278 11234 11133 25 26 9756 MX3X1 $T=1191860 1030330 1 180 $X=1184960 $Y=1030078
X4793 9932 10096 25 9552 26 10189 OAI21X1 $T=1129300 1045090 0 0 $X=1129298 $Y=1044838
X4794 9888 25 74 9914 26 9929 9747 OAI211XL $T=1120560 1310770 0 0 $X=1120558 $Y=1310518
X4795 9952 25 9386 9948 26 9886 9480 OAI211XL $T=1125160 1192690 1 180 $X=1122860 $Y=1192438
X4796 9569 9574 26 9587 25 9659 NOR3BXL $T=1104460 1177930 1 0 $X=1104458 $Y=1173990
X4797 9695 9736 26 9709 25 9906 NOR3BXL $T=1112280 1141030 0 0 $X=1112278 $Y=1140778
X4798 8819 8822 25 8827 8738 26 8818 8870 8953 OAI222XL $T=1057540 1141030 0 0 $X=1057538 $Y=1140778
X4799 8947 8859 25 8677 8940 26 8936 8741 8869 OAI222XL $T=1066740 1148410 1 180 $X=1063060 $Y=1148158
X4800 8943 8931 25 8880 8976 26 8975 9005 9040 OAI222XL $T=1067200 1141030 0 0 $X=1067198 $Y=1140778
X4801 8947 8920 25 8859 8940 26 8936 8677 9066 OAI222XL $T=1068580 1155790 0 0 $X=1068578 $Y=1155538
X4802 8870 9177 25 9141 8931 26 8880 9119 9004 OAI222XL $T=1081000 1141030 1 180 $X=1077320 $Y=1140778
X4803 8943 8947 25 8940 8976 26 8936 9141 9121 OAI222XL $T=1081920 1163170 0 180 $X=1078240 $Y=1159230
X4804 8947 9141 25 9119 8940 26 8936 9353 9521 OAI222XL $T=1094340 1148410 0 0 $X=1094338 $Y=1148158
X4805 9119 8980 25 9353 9243 26 9359 9437 9009 OAI222XL $T=1101700 1141030 1 180 $X=1098020 $Y=1140778
X4806 8951 9432 25 9119 8947 26 8940 9353 9704 OAI222XL $T=1104000 1170550 1 0 $X=1103998 $Y=1166610
X4807 9089 9077 26 9120 9128 25 9145 AOI31X1 $T=1076400 1148410 1 0 $X=1076398 $Y=1144470
.ENDS
***************************************
.SUBCKT ICV_34 3 4 12 13 14 15 16 17 18 19 20 21 22 23 24 42 43 4158
** N=160663 EP=18 IP=47 FDC=0
X0 4 3 12 TIELO $T=746120 749890 0 0 $X=746118 $Y=749638
X1 4 3 15 TIELO $T=747040 749890 0 0 $X=747038 $Y=749638
X2 4 3 16 TIELO $T=747960 749890 0 0 $X=747958 $Y=749638
X3 43 3 4 12941 CLKINVX1 $T=1622420 986050 1 0 $X=1622418 $Y=982110
X4 13 14 4 3 INVX12 $T=746580 749890 1 0 $X=746578 $Y=745950
X5 18 17 4 3 INVX12 $T=750720 749890 1 0 $X=750718 $Y=745950
X6 20 19 4 3 INVX12 $T=752560 757270 1 0 $X=752558 $Y=753330
X7 22 21 4 3 INVX12 $T=754860 749890 1 0 $X=754858 $Y=745950
X8 24 23 4 3 INVX12 $T=759000 749890 1 0 $X=758998 $Y=745950
X9 12941 42 4 3 INVX12 $T=1619200 978670 1 180 $X=1615520 $Y=978418
.ENDS
***************************************
.SUBCKT ICV_35
** N=153840 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_36 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 71 72 73 74 75 76 77 78 79 80 81 82 83 84
+ 85 86 87 88 89 90 91 92 93 94 123
** N=123 EP=91 IP=150 FDC=0
X0 1 41 PDO02CDG $T=251435 0 0 0 $X=255123 $Y=-5002
X1 1 42 PDO02CDG $T=291870 0 0 0 $X=295558 $Y=-5002
X2 1 43 PDO02CDG $T=332305 0 0 0 $X=335993 $Y=-5002
X3 1 44 PDO02CDG $T=372740 0 0 0 $X=376428 $Y=-5002
X4 1 45 PDO02CDG $T=413175 0 0 0 $X=416863 $Y=-5002
X5 2 46 PDO02CDG $T=453610 0 0 0 $X=457298 $Y=-5002
X6 2 47 PDO02CDG $T=494045 0 0 0 $X=497733 $Y=-5002
X7 2 48 PDO02CDG $T=534480 0 0 0 $X=538168 $Y=-5002
X8 2 49 PDO02CDG $T=574915 0 0 0 $X=578603 $Y=-5002
X9 2 50 PDO02CDG $T=615350 0 0 0 $X=619038 $Y=-5002
X10 3 51 PDO02CDG $T=655785 0 0 0 $X=659473 $Y=-5002
X11 3 52 PDO02CDG $T=696220 0 0 0 $X=699908 $Y=-5002
X12 3 53 PDO02CDG $T=736655 0 0 0 $X=740343 $Y=-5002
X13 4 54 PDO02CDG $T=777090 0 0 0 $X=780778 $Y=-5002
X14 5 55 PDO02CDG $T=817525 0 0 0 $X=821213 $Y=-5002
X15 6 56 PDO02CDG $T=857960 0 0 0 $X=861648 $Y=-5002
X16 7 57 PDO02CDG $T=898395 0 0 0 $X=902083 $Y=-5002
X17 8 58 PDO02CDG $T=938830 0 0 0 $X=942518 $Y=-5002
X18 9 59 PDO02CDG $T=979265 0 0 0 $X=982953 $Y=-5002
X19 10 60 PDO02CDG $T=1019700 0 0 0 $X=1023388 $Y=-5002
X20 11 61 PDO02CDG $T=1060135 0 0 0 $X=1063823 $Y=-5002
X21 12 62 PDO02CDG $T=1100565 0 0 0 $X=1104253 $Y=-5002
X22 13 63 PDO02CDG $T=1140995 0 0 0 $X=1144683 $Y=-5002
X23 14 64 PDO02CDG $T=1181425 0 0 0 $X=1185113 $Y=-5002
X24 15 65 PDO02CDG $T=1221855 0 0 0 $X=1225543 $Y=-5002
X25 16 66 PDO02CDG $T=1262285 0 0 0 $X=1265973 $Y=-5002
X26 17 71 PDO02CDG $T=1383575 0 0 0 $X=1387263 $Y=-5002
X27 18 72 PDO02CDG $T=1424005 0 0 0 $X=1427693 $Y=-5002
X28 19 73 PDO02CDG $T=1464435 0 0 0 $X=1468123 $Y=-5002
X29 20 74 PDO02CDG $T=1504865 0 0 0 $X=1508553 $Y=-5002
X30 21 75 PDO02CDG $T=1545300 0 0 0 $X=1548988 $Y=-5002
X31 22 76 PDO02CDG $T=1585735 0 0 0 $X=1589423 $Y=-5002
X32 23 77 PDO02CDG $T=1626170 0 0 0 $X=1629858 $Y=-5002
X33 24 78 PDO02CDG $T=1666605 0 0 0 $X=1670293 $Y=-5002
X34 25 79 PDO02CDG $T=1707040 0 0 0 $X=1710728 $Y=-5002
X35 26 80 PDO02CDG $T=1747475 0 0 0 $X=1751163 $Y=-5002
X36 27 81 PDO02CDG $T=1787910 0 0 0 $X=1791598 $Y=-5002
X37 28 82 PDO02CDG $T=1828345 0 0 0 $X=1832033 $Y=-5002
X38 29 83 PDO02CDG $T=1868780 0 0 0 $X=1872468 $Y=-5002
X39 30 84 PDO02CDG $T=1909215 0 0 0 $X=1912903 $Y=-5002
X40 31 85 PDO02CDG $T=1949650 0 0 0 $X=1953338 $Y=-5002
X41 32 86 PDO02CDG $T=1990085 0 0 0 $X=1993773 $Y=-5002
X42 33 87 PDO02CDG $T=2030520 0 0 0 $X=2034208 $Y=-5002
X43 34 88 PDO02CDG $T=2070955 0 0 0 $X=2074643 $Y=-5002
X44 35 89 PDO02CDG $T=2111390 0 0 0 $X=2115078 $Y=-5002
X45 36 90 PDO02CDG $T=2151825 0 0 0 $X=2155513 $Y=-5002
X46 37 91 PDO02CDG $T=2192260 0 0 0 $X=2195948 $Y=-5002
X47 38 92 PDO02CDG $T=2232695 0 0 0 $X=2236383 $Y=-5002
X48 39 93 PDO02CDG $T=2273130 0 0 0 $X=2276818 $Y=-5002
X49 40 94 PDO02CDG $T=2313565 0 0 0 $X=2317253 $Y=-5002
.ENDS
***************************************
.SUBCKT ICV_37
** N=81 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_38
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_39
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_40 1 2 3 4 5 6 7 11
** N=11 EP=8 IP=15 FDC=0
X0 1 3 PDO02CDG $T=0 2190570 0 270 $X=-5002 $Y=2160850
X1 1 4 PDO02CDG $T=0 2230255 0 270 $X=-5002 $Y=2200535
X2 1 5 PDO02CDG $T=0 2269940 0 270 $X=-5002 $Y=2240220
X3 1 6 PDO02CDG $T=0 2309625 0 270 $X=-5002 $Y=2279905
X4 2 7 PDO02CDG $T=0 2349310 0 270 $X=-5002 $Y=2319590
.ENDS
***************************************
.SUBCKT ICV_41 1 2 3 4 5 6 7 10
** N=10 EP=8 IP=15 FDC=0
X0 2 3 PDO02CDG $T=0 1992145 0 270 $X=-5002 $Y=1962425
X1 2 4 PDO02CDG $T=0 2031830 0 270 $X=-5002 $Y=2002110
X2 2 5 PDO02CDG $T=0 2071515 0 270 $X=-5002 $Y=2041795
X3 1 6 PDO02CDG $T=0 2111200 0 270 $X=-5002 $Y=2081480
X4 1 7 PDO02CDG $T=0 2150885 0 270 $X=-5002 $Y=2121165
.ENDS
***************************************
.SUBCKT ICV_42 1 2 3 4 5 6 7 12
** N=12 EP=8 IP=15 FDC=0
X0 2 3 PDO02CDG $T=0 1793720 0 270 $X=-5002 $Y=1764000
X1 2 4 PDO02CDG $T=0 1833405 0 270 $X=-5002 $Y=1803685
X2 1 5 PDO02CDG $T=0 1873090 0 270 $X=-5002 $Y=1843370
X3 1 6 PDO02CDG $T=0 1912775 0 270 $X=-5002 $Y=1883055
X4 1 7 PDO02CDG $T=0 1952460 0 270 $X=-5002 $Y=1922740
.ENDS
***************************************
.SUBCKT ICV_43 1 2 3 4 5 6 7 9 10 11 12 13 14 15 16 17 18 26
** N=26 EP=18 IP=30 FDC=0
X0 4 9 PDO02CDG $T=0 1396870 0 270 $X=-5002 $Y=1367150
X1 5 10 PDO02CDG $T=0 1436555 0 270 $X=-5002 $Y=1406835
X2 6 11 PDO02CDG $T=0 1476240 0 270 $X=-5002 $Y=1446520
X3 7 12 PDO02CDG $T=0 1515925 0 270 $X=-5002 $Y=1486205
X4 1 13 PDO02CDG $T=0 1555610 0 270 $X=-5002 $Y=1525890
X5 2 14 PDO02CDG $T=0 1595295 0 270 $X=-5002 $Y=1565575
X6 3 15 PDO02CDG $T=0 1634980 0 270 $X=-5002 $Y=1605260
X7 3 16 PDO02CDG $T=0 1674665 0 270 $X=-5002 $Y=1644945
X8 3 17 PDO02CDG $T=0 1714350 0 270 $X=-5002 $Y=1684630
X9 3 18 PDO02CDG $T=0 1754035 0 270 $X=-5002 $Y=1724315
.ENDS
***************************************
.SUBCKT ICV_44 1 2 3 4 5 6 7 8 9 10 11 12 13 14 22
** N=24 EP=15 IP=21 FDC=0
X0 1 8 PDO02CDG $T=0 1039705 0 270 $X=-5002 $Y=1009985
X1 2 9 PDO02CDG $T=0 1079390 0 270 $X=-5002 $Y=1049670
X2 3 10 PDO02CDG $T=0 1119075 0 270 $X=-5002 $Y=1089355
X3 4 11 PDO02CDG $T=0 1158760 0 270 $X=-5002 $Y=1129040
X4 5 12 PDO02CDG $T=0 1198445 0 270 $X=-5002 $Y=1168725
X5 6 13 PDO02CDG $T=0 1238130 0 270 $X=-5002 $Y=1208410
X6 7 14 PDO02CDG $T=0 1277815 0 270 $X=-5002 $Y=1248095
.ENDS
***************************************
.SUBCKT ICV_45 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 23
** N=23 EP=19 IP=27 FDC=0
X0 1 10 PDO02CDG $T=0 682540 0 270 $X=-5002 $Y=652820
X1 2 11 PDO02CDG $T=0 722225 0 270 $X=-5002 $Y=692505
X2 3 12 PDO02CDG $T=0 761910 0 270 $X=-5002 $Y=732190
X3 4 13 PDO02CDG $T=0 801595 0 270 $X=-5002 $Y=771875
X4 5 14 PDO02CDG $T=0 841280 0 270 $X=-5002 $Y=811560
X5 6 15 PDO02CDG $T=0 880965 0 270 $X=-5002 $Y=851245
X6 7 16 PDO02CDG $T=0 920650 0 270 $X=-5002 $Y=890930
X7 8 17 PDO02CDG $T=0 960335 0 270 $X=-5002 $Y=930615
X8 9 18 PDO02CDG $T=0 1000020 0 270 $X=-5002 $Y=970300
.ENDS
***************************************
.SUBCKT ICV_46 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 26
** N=26 EP=21 IP=30 FDC=0
X0 1 11 PDO02CDG $T=0 285690 0 270 $X=-5002 $Y=255970
X1 2 12 PDO02CDG $T=0 325375 0 270 $X=-5002 $Y=295655
X2 3 13 PDO02CDG $T=0 365060 0 270 $X=-5002 $Y=335340
X3 4 14 PDO02CDG $T=0 404745 0 270 $X=-5002 $Y=375025
X4 5 15 PDO02CDG $T=0 444430 0 270 $X=-5002 $Y=414710
X5 6 16 PDO02CDG $T=0 484115 0 270 $X=-5002 $Y=454395
X6 7 17 PDO02CDG $T=0 523800 0 270 $X=-5002 $Y=494080
X7 8 18 PDO02CDG $T=0 563485 0 270 $X=-5002 $Y=533765
X8 9 19 PDO02CDG $T=0 603170 0 270 $X=-5002 $Y=573450
X9 10 20 PDO02CDG $T=0 642855 0 270 $X=-5002 $Y=613135
.ENDS
***************************************
.SUBCKT ICV_47
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_48
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_49
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_50
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_51
** N=10 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_52
** N=12 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_53
** N=11 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_54
** N=20 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_55
** N=17 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_56
** N=18 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_57
** N=17 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_58
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_59
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CHIP VDD VSS DCACHE_rdata[13] DCACHE_rdata[16] DCACHE_rdata[15] DCACHE_rdata[14] DCACHE_rdata[17] DCACHE_rdata[18] DCACHE_rdata[22] DCACHE_rdata[21] DCACHE_rdata[20] DCACHE_rdata[19] DCACHE_rdata[23] DCACHE_rdata[26] DCACHE_rdata[25] DCACHE_rdata[24] DCACHE_rdata[27] DCACHE_rdata[28] test_so DCACHE_wen
+ DCACHE_ren ICACHE_wen ICACHE_ren DCACHE_rdata[31] DCACHE_rdata[30] DCACHE_rdata[29] ICACHE_addr[7] ICACHE_addr[6] ICACHE_addr[5] ICACHE_addr[4] ICACHE_addr[3] ICACHE_addr[2] ICACHE_addr[1] ICACHE_addr[0] ICACHE_addr[8] ICACHE_addr[16] ICACHE_addr[15] ICACHE_addr[14] ICACHE_addr[13] ICACHE_addr[12]
+ ICACHE_addr[11] ICACHE_addr[10] ICACHE_addr[9] ICACHE_addr[17] ICACHE_addr[26] ICACHE_addr[25] ICACHE_addr[24] ICACHE_addr[23] ICACHE_addr[22] ICACHE_addr[21] ICACHE_addr[20] ICACHE_addr[19] ICACHE_addr[18] DCACHE_rdata[12] ICACHE_addr[27] ICACHE_rdata[0] ICACHE_rdata[1] ICACHE_rdata[2] ICACHE_rdata[3] ICACHE_rdata[4]
+ ICACHE_rdata[5] ICACHE_rdata[6] ICACHE_rdata[7] ICACHE_rdata[8] ICACHE_rdata[9] ICACHE_rdata[10] ICACHE_rdata[11] ICACHE_rdata[12] ICACHE_rdata[13] ICACHE_rdata[14] ICACHE_rdata[15] ICACHE_rdata[16] ICACHE_rdata[17] ICACHE_rdata[18] ICACHE_rdata[19] ICACHE_rdata[20] ICACHE_rdata[21] ICACHE_rdata[22] ICACHE_rdata[23] ICACHE_rdata[24]
+ ICACHE_rdata[25] ICACHE_rdata[26] ICACHE_rdata[27] ICACHE_rdata[28] ICACHE_rdata[29] ICACHE_rdata[30] ICACHE_rdata[31] clk rst ICACHE_stall DCACHE_stall test_si test_se DCACHE_rdata[0] DCACHE_rdata[1] DCACHE_rdata[2] DCACHE_rdata[3] DCACHE_rdata[4] DCACHE_rdata[5] DCACHE_rdata[6]
+ DCACHE_rdata[7] DCACHE_rdata[8] DCACHE_rdata[9] DCACHE_rdata[10] DCACHE_rdata[11] ICACHE_wdata[12] ICACHE_wdata[11] ICACHE_wdata[10] ICACHE_wdata[9] ICACHE_wdata[8] ICACHE_wdata[7] ICACHE_wdata[6] ICACHE_wdata[5] ICACHE_wdata[4] ICACHE_wdata[3] ICACHE_wdata[2] ICACHE_wdata[1] ICACHE_wdata[0] DCACHE_addr[31] DCACHE_addr[30]
+ DCACHE_addr[29] DCACHE_addr[28] DCACHE_addr[27] DCACHE_addr[26] DCACHE_addr[25] DCACHE_addr[24] DCACHE_addr[23] DCACHE_addr[22] DCACHE_addr[21] DCACHE_addr[20] DCACHE_addr[19] DCACHE_addr[18] DCACHE_addr[17] DCACHE_addr[16] DCACHE_addr[15] DCACHE_addr[14] DCACHE_addr[13] DCACHE_addr[12] DCACHE_addr[11] DCACHE_addr[10]
+ DCACHE_addr[9] DCACHE_addr[8] DCACHE_addr[7] DCACHE_addr[6] DCACHE_addr[5] DCACHE_addr[4] DCACHE_addr[3] DCACHE_addr[2] DCACHE_addr[1] DCACHE_addr[0] ICACHE_addr[31] ICACHE_addr[30] ICACHE_addr[29] ICACHE_addr[28] ICACHE_wdata[17] ICACHE_wdata[16] ICACHE_wdata[15] ICACHE_wdata[14] ICACHE_wdata[13] ICACHE_wdata[22]
+ ICACHE_wdata[21] ICACHE_wdata[20] ICACHE_wdata[19] ICACHE_wdata[18] ICACHE_wdata[27] ICACHE_wdata[26] ICACHE_wdata[25] ICACHE_wdata[24] ICACHE_wdata[23] DCACHE_wdata[5] DCACHE_wdata[4] DCACHE_wdata[3] DCACHE_wdata[2] DCACHE_wdata[1] DCACHE_wdata[0] ICACHE_wdata[31] ICACHE_wdata[30] ICACHE_wdata[29] ICACHE_wdata[28] DCACHE_wdata[12]
+ DCACHE_wdata[11] DCACHE_wdata[10] DCACHE_wdata[9] DCACHE_wdata[8] DCACHE_wdata[7] DCACHE_wdata[6] DCACHE_wdata[21] DCACHE_wdata[20] DCACHE_wdata[19] DCACHE_wdata[18] DCACHE_wdata[17] DCACHE_wdata[16] DCACHE_wdata[15] DCACHE_wdata[14] DCACHE_wdata[13] DCACHE_wdata[31] DCACHE_wdata[30] DCACHE_wdata[29] DCACHE_wdata[28] DCACHE_wdata[27]
+ DCACHE_wdata[26] DCACHE_wdata[25] DCACHE_wdata[24] DCACHE_wdata[23] DCACHE_wdata[22]
** N=12196 EP=205 IP=24886 FDC=0
X13 3279 3280 4135 4133 4134 DCACHE_rdata[17] DCACHE_rdata[16] DCACHE_rdata[15] DCACHE_rdata[14] DCACHE_rdata[13] 12196 ICV_14 $T=0 0 0 0 $X=2354000 $Y=2160800
X14 4852 3281 1159 3282 3283 DCACHE_rdata[22] DCACHE_rdata[21] DCACHE_rdata[20] DCACHE_rdata[19] DCACHE_rdata[18] 12196 ICV_15 $T=0 0 0 0 $X=2354000 $Y=1962400
X15 1499 1377 1374 1376 1497 DCACHE_rdata[27] DCACHE_rdata[26] DCACHE_rdata[25] DCACHE_rdata[24] DCACHE_rdata[23] 12196 ICV_16 $T=0 0 0 0 $X=2354000 $Y=1763998
X16 1 2 3287 3288 3289 9296 3284 3285 3286 test_so DCACHE_wen DCACHE_ren ICACHE_wen ICACHE_ren DCACHE_rdata[31] DCACHE_rdata[30] DCACHE_rdata[29] DCACHE_rdata[28] 12196 ICV_17 $T=0 0 0 0 $X=2354000 $Y=1351600
X17 8432 8431 8427 8229 8426 5522 8271 8434 ICACHE_addr[7] ICACHE_addr[6] ICACHE_addr[5] ICACHE_addr[4] ICACHE_addr[3] ICACHE_addr[2] ICACHE_addr[1] ICACHE_addr[0] 12196 ICV_18 $T=0 0 0 0 $X=2354000 $Y=1008393
X18 3 8433 1853 5126 8272 8430 5153 8429 8428 ICACHE_addr[16] ICACHE_addr[15] ICACHE_addr[14] ICACHE_addr[13] ICACHE_addr[12] ICACHE_addr[11] ICACHE_addr[10] ICACHE_addr[9] ICACHE_addr[8] 12196 ICV_19 $T=0 0 0 0 $X=2354000 $Y=639200
X19 2383 5762 9296 1814 8621 8592 8259 8784 8247 2391 ICACHE_addr[26] ICACHE_addr[25] ICACHE_addr[24] ICACHE_addr[23] ICACHE_addr[22] ICACHE_addr[21] ICACHE_addr[20] ICACHE_addr[19] ICACHE_addr[18] ICACHE_addr[17]
+ 12196
+ ICV_20 $T=0 0 0 0 $X=2354000 $Y=246000
X23 3854 484 485 486 487 488 489 490 3855 3856 3857 3858 491 3859 3860 3861 608 492 493 494
+ 495 3862 3863 7101 496 497 3864 498 3865 499 500 501 3866 502 503 504 505 3867 506 507
+ 508 509 510 511 512 513 514 515 516 517 518 ICACHE_rdata[0] ICACHE_rdata[1] ICACHE_rdata[2] ICACHE_rdata[3] ICACHE_rdata[4] ICACHE_rdata[5] ICACHE_rdata[6] ICACHE_rdata[7] ICACHE_rdata[8]
+ ICACHE_rdata[9] ICACHE_rdata[10] ICACHE_rdata[11] ICACHE_rdata[12] ICACHE_rdata[13] ICACHE_rdata[14] ICACHE_rdata[15] ICACHE_rdata[16] ICACHE_rdata[17] ICACHE_rdata[18] ICACHE_rdata[19] ICACHE_rdata[20] ICACHE_rdata[21] ICACHE_rdata[22] ICACHE_rdata[23] ICACHE_rdata[24] ICACHE_rdata[25] ICACHE_rdata[26] ICACHE_rdata[27] ICACHE_rdata[28]
+ ICACHE_rdata[29] ICACHE_rdata[30] ICACHE_rdata[31] clk rst ICACHE_stall DCACHE_stall test_si test_se DCACHE_rdata[0] DCACHE_rdata[1] DCACHE_rdata[2] DCACHE_rdata[3] DCACHE_rdata[4] DCACHE_rdata[5] DCACHE_rdata[6] DCACHE_rdata[7] DCACHE_rdata[8] DCACHE_rdata[9] DCACHE_rdata[10]
+ DCACHE_rdata[11] DCACHE_rdata[12] 12196
+ ICV_24 $T=0 0 0 0 $X=246000 $Y=2354000
X26 VSS VDD 262 4 5 4723 3866 1381 503 504 12196 ICV_27 $T=0 0 0 0 $X=246000 $Y=1764000
X27 284 VSS VDD 1591 282 283 1627 1705 1661 5029 1666 1667 5066 493 1668 5020 1670 494 1671 492
+ 5028 5024 1672 1673 5021 608 1669 1674 5035 495 1677 1676 5050 3860 1663 5030 1678 5033 1679 1680
+ 3862 3858 484 5045 3859 1708 3861 5032 3857 5031 1683 5037 1685 1686 1699 491 5036 5095 1688 5053
+ 1689 1949 1691 5039 7101 487 1714 5042 5043 5060 5038 1695 486 5040 5046 1703 1702 488 1706 5151
+ 1704 1707 5051 5055 8250 489 5082 1710 485 1662 5072 5067 5047 1724 3856 1716 5065 1717 1719 490
+ 5088 3854 1722 5070 8263 1733 5080 5075 1723 3863 496 1712 5077 1725 5073 1730 1726 5068 5083 1728
+ 3855 1729 497 1731 5081 5089 5058 5094 1736 5086 1737 5091 1727 1740 1777 5195 5092 8784 8259 1741
+ 1742 1743 3865 3864 5096 5090 8208 498 1747 8206 1748 499 8433 5108 5101 5117 5098 1745 500 5099
+ 501 1749 5113 1750 1853 5119 1812 1751 8221 5102 1753 1752 1759 1755 8272 1756 1758 5109 5126 3
+ 8213 1761 5115 1762 1764 8430 5111 6953 505 1766 5120 5123 1767 5125 8429 2400 5093 5129 5127 5137
+ 1774 1772 5136 8215 1775 5132 1830 1776 8214 1765 2526 1778 1771 5159 5134 1780 5135 1781 8434 5140
+ 8222 5139 5153 1783 1773 5142 1794 5144 1782 5143 1787 5145 5133 1789 1785 1788 1790 5158 5147 1792
+ 1793 2518 1795 5152 1796 1805 8229 8234 1797 8271 5150 5149 1808 5173 5176 5160 5166 1828 8432 1800
+ 1802 5232 1804 8426 5231 1807 1843 8428 5165 8247 1801 1815 6957 5182 1806 8245 5141 5161 6954 1809
+ 5235 5171 5245 1823 1811 5169 5167 5271 5162 5239 5163 5172 6956 1954 1814 5184 1816 8236 1831 5187
+ 1819 5179 5177 1822 5189 4723 1820 1825 1826 5185 1829 5298 1952 5180 5196 5188 1967 5313 1833 5236
+ 5312 5194 8275 5191 1893 1847 1835 1836 5308 5280 5242 1890 1845 8274 5335 8268 5285 1972 1837 8427
+ 1838 5330 8244 1860 5217 1842 1841 8431 5199 5197 8249 5219 1846 1844 1848 5203 5202 8246 5218 8253
+ 5320 5224 5200 5315 1849 1850 5156 8251 5221 1851 5213 5121 5205 3725 5292 5283 5309 5264 5268 5223
+ 5253 5248 1857 5130 5230 5148 5346 5215 1863 1861 1855 5222 5124 5128 5210 8248 1862 5104 5174 5154
+ 1866 5107 8220 5118 8252 5267 1865 1871 1878 1869 5211 5229 5216 5522 5228 5226 1872 1873 1978 5238
+ 1874 8258 1875 5227 1903 5251 1876 5241 1877 1883 1895 1885 1879 1881 1889 5225 1888 1887 1897 1886
+ 3683 5249 1891 5252 1892 5246 5282 1909 1905 1964 5254 1899 5290 1900 5257 5261 5269 5263 1896 1930
+ 1906 8267 5293 5256 1931 5262 5275 5270 5302 1914 1922 5279 5289 5300 5281 1911 1910 1915 1916 5304
+ 1917 1945 5284 1918 1919 5277 5286 1923 1924 5311 1926 1934 1927 1973 1944 1929 5307 5297 5288 1933
+ 5295 1953 5314 1942 1955 1959 8278 5301 1943 1936 1950 1938 1937 1939 5332 1940 5316 1948 1951 8273
+ 5321 1976 1960 8283 5317 1961 8285 1957 5319 1979 1962 5322 8282 5324 5328 1966 5325 5326 5323 5329
+ 1971 8284 1963 1968 1969 3867 5333 5331 1980 1981 5336 1984 1965 2001 5327 1989 1983 5338 2008 5343
+ 1992 1985 2391 5351 1990 5345 1991 5344 1997 1996 1998 2007 5359 3287 1999 5349 5353 3289 2 3288
+ 5354 2002 2010 2004 1374 2006 2005 2009 517 512 516 1376 2011 2014 1995 1993 2013 2012 515 511
+ 513 502 2015 510 1381 3284 1 3285 3286 12196
+ ICV_30 $T=0 0 0 0 $X=246000 $Y=1351110
X28 VSS VDD 2257 1672 1668 5029 1661 1662 1663 1669 2167 1667 1591 2258 1670 2265 5020 1666 5021 1671
+ 5624 1627 2259 1673 1674 5058 5673 5028 5024 1676 5668 5674 1677 2256 1705 1678 1679 1680 2260 5030
+ 3797 5036 1683 1708 1686 5633 1699 5031 2169 5051 5661 1685 5035 5033 5032 2303 5039 1695 5037 1688
+ 5066 1689 5675 5043 5038 1949 1706 5040 1691 2168 5047 5042 3742 5046 1788 3173 3741 1707 1714 1704
+ 1702 1703 5050 3743 8583 1722 5691 5055 5524 1710 5045 1712 5702 5095 3744 1717 1716 5065 7019 8626
+ 5067 5077 5525 7022 5068 3748 7017 3746 3745 1723 7021 7018 5093 1724 5727 5073 1725 1726 5737 1727
+ 5078 1728 1805 1729 5080 5072 5081 7020 1730 1734 5084 1731 3747 1736 1765 5070 5086 1773 5075 5088
+ 5092 1743 5090 1749 1777 1740 5091 1741 1737 8592 3697 5085 5845 5096 8206 1745 1747 5098 1748 5053
+ 1869 5107 1751 1742 5099 5101 5060 1719 1750 5104 8208 1752 5113 5102 5111 1753 1776 1755 1767 1761
+ 1756 1733 1759 5133 1758 1766 8214 1771 5752 1762 5118 5119 5132 6957 5162 5142 5083 1764 5121 5128
+ 5127 5124 2492 5141 5151 1828 2482 1780 1772 5130 2474 5115 8215 1778 5135 5134 5798 2462 1830 5137
+ 1787 5120 1781 1782 5140 5136 1775 8245 8220 5143 5139 1783 1785 2510 5145 5149 5174 5245 1789 2442
+ 5125 5147 1795 1774 1790 8222 5154 5148 5150 5156 1793 5345 1792 1794 8650 2417 1954 1797 1796 2434
+ 5232 1815 5163 8621 6263 6953 5089 5160 1804 5094 1802 6954 1800 5173 5161 2407 1808 8221 1801 5176
+ 5169 5179 5271 5751 2425 1819 5108 5172 5167 5166 5082 5159 5239 1807 5180 5182 2402 5713 5762 1809
+ 2001 5129 5171 1811 1812 5343 8234 1820 5117 5191 1825 5187 5189 5177 5196 1831 2383 8246 1829 5197
+ 1822 1823 5200 5184 1826 8251 5185 1890 1833 5238 1997 5188 8213 1841 5217 1951 8273 5203 1835 1893
+ 1952 5280 1836 5335 8249 5194 5285 1985 5314 5298 5219 5312 5236 8253 5195 1816 8258 1838 1837 1845
+ 8268 5242 8244 5224 5321 1846 1842 1843 5199 1844 2008 5202 1847 5320 8248 1848 5221 1849 1851 1915
+ 1850 5230 1862 5210 5225 5264 8252 5309 5292 3725 5313 5268 5223 5218 5205 1877 1857 5248 8250 5211
+ 1855 1861 5227 1860 5267 5222 5213 5109 5229 1814 5215 1863 1866 5216 1865 5165 5123 1873 1874 1913
+ 1875 1871 1872 5226 1876 1886 5228 1883 5246 5253 1879 5231 5158 5315 1889 1878 5235 1881 5241 5144
+ 1891 1885 1903 1887 5254 3683 1888 1892 1899 1897 5256 1896 1895 5261 8263 5249 1900 5257 5252 5251
+ 1972 5282 5263 1922 1906 6956 5269 4723 5262 1909 8267 5275 1905 1910 5279 1930 1914 1911 5289 5270
+ 5277 1916 1917 1919 1918 5152 5304 1931 5281 5284 5288 5316 5286 1927 5300 1923 5311 1926 5283 1924
+ 1929 5295 5290 1933 5297 1942 1934 1936 1944 5301 5322 1950 5293 5302 2518 2526 1937 1938 1939 1943
+ 1940 5332 1978 1953 1945 5330 8274 1948 8275 5308 5307 8278 1955 5317 5324 1957 1965 1963 1960 8285
+ 1961 5319 1979 1962 1964 5323 8282 5329 1966 5325 5338 1971 1967 5327 1969 8283 1968 1980 5331 1973
+ 8284 1984 1959 5333 1976 5326 5328 1981 5336 1983 5351 2391 1989 8236 1990 1992 5344 1993 1991 2004
+ 1996 1995 5349 1998 1999 2010 5354 5353 2011 2002 5346 3282 3 3279 5359 2005 1499 2009 4133 1159
+ 2007 2015 2006 3281 1377 2012 3283 4135 2014 3280 508 2013 4134 4852 518 1497 507 514 509 506
+ 9296 12196
+ ICV_33 $T=0 0 0 0 $X=246000 $Y=1008400
X29 VSS VDD 2695 2256 376 2694 2693 372 2257 373 2258 375 2259 374 2260 2400 1806 12196 ICV_34 $T=0 0 0 0 $X=246000 $Y=639200
X31 2695 2694 2693 2265 5624 5633 8583 5674 5673 2303 5661 5668 5675 3173 5691 5702 8626 5727 5737 6263
+ 8650 5751 2402 2407 2417 2425 2434 2442 5798 2462 2474 2482 2492 5752 5845 5713 2510 2518 2526 2400
+ ICACHE_wdata[12] ICACHE_wdata[11] ICACHE_wdata[10] ICACHE_wdata[9] ICACHE_wdata[8] ICACHE_wdata[7] ICACHE_wdata[6] ICACHE_wdata[5] ICACHE_wdata[4] ICACHE_wdata[3] ICACHE_wdata[2] ICACHE_wdata[1] ICACHE_wdata[0] DCACHE_addr[31] DCACHE_addr[30] DCACHE_addr[29] DCACHE_addr[28] DCACHE_addr[27] DCACHE_addr[26] DCACHE_addr[25]
+ DCACHE_addr[24] DCACHE_addr[23] DCACHE_addr[22] DCACHE_addr[21] DCACHE_addr[20] DCACHE_addr[19] DCACHE_addr[18] DCACHE_addr[17] DCACHE_addr[16] DCACHE_addr[15] DCACHE_addr[14] DCACHE_addr[13] DCACHE_addr[12] DCACHE_addr[11] DCACHE_addr[10] DCACHE_addr[9] DCACHE_addr[8] DCACHE_addr[7] DCACHE_addr[6] DCACHE_addr[5]
+ DCACHE_addr[4] DCACHE_addr[3] DCACHE_addr[2] DCACHE_addr[1] DCACHE_addr[0] ICACHE_addr[31] ICACHE_addr[30] ICACHE_addr[29] ICACHE_addr[28] ICACHE_addr[27] 12196
+ ICV_36 $T=0 0 0 0 $X=246000 $Y=-5002
X35 4 5 ICACHE_wdata[17] ICACHE_wdata[16] ICACHE_wdata[15] ICACHE_wdata[14] ICACHE_wdata[13] 12196 ICV_40 $T=0 0 0 0 $X=-5002 $Y=2160800
X36 4 262 ICACHE_wdata[22] ICACHE_wdata[21] ICACHE_wdata[20] ICACHE_wdata[19] ICACHE_wdata[18] 12196 ICV_41 $T=0 0 0 0 $X=-5002 $Y=1962400
X37 262 284 ICACHE_wdata[27] ICACHE_wdata[26] ICACHE_wdata[25] ICACHE_wdata[24] ICACHE_wdata[23] 12196 ICV_42 $T=0 0 0 0 $X=-5002 $Y=1764000
X38 282 283 284 1734 5078 5084 5085 DCACHE_wdata[5] DCACHE_wdata[4] DCACHE_wdata[3] DCACHE_wdata[2] DCACHE_wdata[1] DCACHE_wdata[0] ICACHE_wdata[31] ICACHE_wdata[30] ICACHE_wdata[29] ICACHE_wdata[28] 12196 ICV_43 $T=0 0 0 0 $X=-5002 $Y=1351600
X39 7017 7018 7019 3697 7020 7021 7022 DCACHE_wdata[12] DCACHE_wdata[11] DCACHE_wdata[10] DCACHE_wdata[9] DCACHE_wdata[8] DCACHE_wdata[7] DCACHE_wdata[6] 12196 ICV_44 $T=0 0 0 0 $X=-5002 $Y=1008400
X40 3741 3742 3743 3744 5525 3745 3746 3747 3748 DCACHE_wdata[21] DCACHE_wdata[20] DCACHE_wdata[19] DCACHE_wdata[18] DCACHE_wdata[17] DCACHE_wdata[16] DCACHE_wdata[15] DCACHE_wdata[14] DCACHE_wdata[13] 12196 ICV_45 $T=0 0 0 0 $X=-5002 $Y=639200
X41 372 373 374 375 376 2167 5524 2168 2169 3797 DCACHE_wdata[31] DCACHE_wdata[30] DCACHE_wdata[29] DCACHE_wdata[28] DCACHE_wdata[27] DCACHE_wdata[26] DCACHE_wdata[25] DCACHE_wdata[24] DCACHE_wdata[23] DCACHE_wdata[22]
+ 12196
+ ICV_46 $T=0 0 0 0 $X=-5002 $Y=246000
.ENDS
***************************************
