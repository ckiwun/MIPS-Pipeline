   module RF2SH64x16 ( 
   	QA,
	DB,
	CLKB,
	CLKA,
	CENB,
	CENA,
	AB,		
	AA);
	
	output	[15:0]	QA;
	input	[15:0]	DB;
	input	CLKB;
	input	CLKA;
	input	CENB;
	input	CENA;
	input	[5:0]	AB;		
	input	[5:0]	AA;
	
	endmodule
	
	
	
